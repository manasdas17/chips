--+============================================================================+
--|                   *** SVGA CHARACTER DISPLAY ***                           |
--+============================================================================+
--| Filename         :svga_core.vhd                                            |
--| Project          :SVGA CHARATER DISPLAY                                    |
--| Version          :0.1                                                      |
--| Author           :Jonathan P Dawson                                        |
--| Created Date     :2005-12-18                                               |
--+============================================================================+
--| Description      :A Python Streams compatible VGA core.                    |
--|                   The core is implemented using BLOCK RAMs to create       |
--|                   character maped graphics. An SVGA (800x600 75hz) display |
--|                   is generated consisting of 100x75 characters of 8x8      |
--|                   pixels each. Each caracter is set to an 8-bit value. At  |
--|                   present ASCII glyphs have been generated.                |
--+============================================================================+
--| Dependencies     :Standard Libraries                                       |
--+============================================================================+
--| Revision History :                                                         |
--|                                                                            |
--| Date :2005-12-18                                                          |
--| Author :Jonathan P Dawson                                                  |
--| Modification: Created File                                                 |
--|                                                                            |
--| Date :2010-12-21                                                           |
--| Author :Jonathan P Dawson                                                  |
--| Modification: Modified for incorporation into Python Streams               |
--|                                                                            |
--+============================================================================+
--| Copyright (C) Jonathan P Dawson 2005                                       |
--+============================================================================+

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity VIDEO_TIME_GEN is
  port ( 
  CLK                    : in  Std_logic;
  RST                    : in  Std_logic;
  CHARADDR               : out Std_logic_vector(12 downto 0);
  PIXROW                 : out Std_logic_vector(2 downto 0);
  PIXCOL                 : out Std_logic_vector(2 downto 0);
  HSYNCH                 : out Std_logic;
  VSYNCH                 : out Std_logic;
  BLANK                  : out Std_logic);
end VIDEO_TIME_GEN;

architecture RTL of VIDEO_TIME_GEN is
  
  signal PIX_ROW_ADDRESS : Unsigned(2 downto 0);
  signal PIX_COL_ADDRESS : Unsigned(2 downto 0);
  signal ROW_ADDRESS     : Unsigned(12 downto 0);
  signal COL_ADDRESS     : Unsigned(6 downto 0);
  
  signal VTIMER          : Unsigned(9 downto 0);
  signal HTIMER          : Unsigned(10 downto 0);
  signal VTIMER_EN       : Std_logic;
  signal VBLANK          : Std_logic;
  signal HBLANK          : Std_logic;
  signal INTVSYNCH       : Std_logic;
  signal INTHSYNCH       : Std_logic;
  
  constant HSYNCHTIME    : Integer := 120;
  constant HACTIVETIME   : Integer := 800;
  constant FPORCHTIME    : Integer := 64;
  constant BPORCHTIME    : Integer := 56;
  
  constant VSYNCHTIME    : Integer := 6;
  constant VACTIVETIME   : Integer := 600;
  constant VFPORCHTIME   : Integer := 35;
  constant VBPORCHTIME   : Integer := 21;
  
begin
  
  process(CLK, RST)
  begin
    if RST = '1' then
      PIX_COL_ADDRESS <= (others => '0');
      PIX_ROW_ADDRESS <= (others => '0');
      COL_ADDRESS     <= (others => '0');
      ROW_ADDRESS     <= (others => '0');
    elsif Rising_edge(CLK) then
      if VBLANK = '0' and HBLANK = '0' then
        if PIX_COL_ADDRESS = To_unsigned(7, 3) then
          PIX_COL_ADDRESS <= (others => '0');
          if COL_ADDRESS = To_unsigned(99, 7) then
            COL_ADDRESS <= (others => '0');
            if PIX_ROW_ADDRESS = To_unsigned(7, 3) then
              PIX_ROW_ADDRESS <= (others => '0');
              if ROW_ADDRESS = To_unsigned(7400, 13) then
                ROW_ADDRESS <= (others => '0');
              else
                ROW_ADDRESS <= ROW_ADDRESS + 100;
              end if;
            else
              PIX_ROW_ADDRESS <= PIX_ROW_ADDRESS + 1;
            end if;
          else
            COL_ADDRESS <= COL_ADDRESS + 1;
          end if;
        else
          PIX_COL_ADDRESS <= PIX_COL_ADDRESS +1;
        end if;
      end if;
    end if;
  end process;
  
  process(CLK, RST)
  begin
    if RST = '1' then
      VTIMER <= (others => '0');
      INTVSYNCH <= '0';
      VBLANK <= '1';
    elsif Rising_edge(CLK) then
      if VTIMER_EN = '1' then
        VTIMER <= VTIMER + 1;
        
        if VTIMER = To_unsigned(VSYNCHTIME, 10) then
          INTVSYNCH <= '1';
        end if;
        
        if VTIMER = To_unsigned(VSYNCHTIME 
          + VFPORCHTIME, 10) then
          VBLANK   <= '0';
        end if;
        
        if VTIMER = To_unsigned(VSYNCHTIME 
          + VFPORCHTIME 
          + VACTIVETIME, 10) then
          VBLANK   <= '1';
        end if;
        
        if VTIMER = To_unsigned(VSYNCHTIME 
          + VFPORCHTIME 
          + VACTIVETIME 
          + VBPORCHTIME, 10) then          
          INTVSYNCH <= '0';
          VTIMER <= (others => '0');
        end if;
      end if;
    end if;
  end process;
  
  process(CLK, RST)
  begin         
    if RST = '1' then
      HTIMER     <= (others => '0');
      INTHSYNCH   <= '0';
      HBLANK   <= '1';
      VTIMER_EN  <= '1';
    elsif Rising_edge(CLK) then
      HTIMER <= HTIMER + 1;
      VTIMER_EN <= '0';
      
      if HTIMER = To_unsigned(HSYNCHTIME, 11) then      
        INTHSYNCH <= '1';
      end if;
      
      if HTIMER = To_unsigned(HSYNCHTIME 
        + FPORCHTIME, 11) then
        HBLANK <= '0';
      end if;
      
      if HTIMER = To_unsigned(HSYNCHTIME 
        + FPORCHTIME 
        + HACTIVETIME, 11) then
        HBLANK <= '1';
      end if;
      
      if HTIMER = To_unsigned(HSYNCHTIME 
        + FPORCHTIME 
        + HACTIVETIME 
        + BPORCHTIME, 11) then          
        INTHSYNCH <= '0';
        VTIMER_EN <= '1';
        HTIMER <= (others => '0');          
      end if;
    end if;              
  end process;
  
  HSYNCH <= INTHSYNCH;
  VSYNCH <= INTVSYNCH;
  BLANK <= HBLANK or VBLANK;
  
  CHARADDR <= Std_logic_vector(ROW_ADDRESS + COL_ADDRESS);
  PIXCOL   <= Std_logic_vector(PIX_COL_ADDRESS);
  PIXROW   <= Std_logic_vector(PIX_ROW_ADDRESS);
  
  
end RTL;

library IEEE;
use Ieee.std_logic_1164.all;
use Ieee.numeric_std.all;

entity CHARACTER_SVGA is
  port ( 

  CLK         : in  Std_logic;
  RST         : in  Std_logic;
  TIMER_1us   : in  Std_logic;
  TIMER_10us  : in  Std_logic;
  TIMER_100us : in  Std_logic;
  TIMER_1ms   : in  Std_logic;

  --Python Streams Interface
  DATA        : in  Std_logic_vector(7 downto 0);
  DATA_STB    : in  Std_logic;
  DATA_ACK    : out Std_logic;
  
  --VGA interface
  R           : out Std_logic;
  G           : out Std_logic;
  B           : out Std_logic;
  HSYNCH      : out Std_logic;
  VSYNCH      : out Std_logic
  );
end CHARACTER_SVGA;

architecture RTL of CHARACTER_SVGA is

  type PIX_ARRAY_TYPE  is array (0 to 2047) of Std_logic_vector(7 downto 0);  
  
  constant PIXARRAY : PIX_ARRAY_TYPE := (
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --0d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --1d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --2d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --3d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --4d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --5d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --6d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --7d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --8d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --9d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --10d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --11d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --12d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --13d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --14d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --15d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --16d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --17d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --18d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --19d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --20d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --21d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --22d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --23d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --24d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --25d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --26d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --27d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --28d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --29d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --30d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --31d
  
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --space
  "00001000","00001000","00001000","00001000","00000000","00001000","00000000","00000000", --!
  "00010100","00010100","00000000","00000000","00000000","00000000","00000000","00000000", --"
  "00000000","00010100","00111110","00010100","00111110","00010100","00000000","00000000", --#
  "00001000","00111100","00001010","00011100","00101000","00011110","00001000","00000000", --$
  "10001110","01001010","00101110","00010000","11101000","10100100","11100010","00000000", --%
  "00001100","00010010","00010010","00001100","00110010","00010010","01101100","00000000", ----'
  "00001000","00001000","00000000","00000000","00000000","00000000","00000000","00000000", --(
  "00001000","00000100","00000010","00000010","00000010","00000100","00001000","00000000", --)
  "00001000","00010000","00100000","00100000","00100000","00010000","00001000","00000000", --*
  "00001000","00111110","00010100","00100010","00000000","00000000","00000000","00000000", --+
  "00010000","00010000","00010000","11111110","00010000","00010000","00010000","00000000", --,
  "00000000","00000000","00000000","00000000","00000000","00001000","00001000","00000000", ---
  "00000000","00000000","00000000","00111110","00000000","00000000","00000000","00000000", --.
  "00000000","00000000","00000000","00000000","00000000","00001000","00000000","00000000", --/
  "01000000","00100000","00010000","00001000","00000100","00000010","00000000","00000000", --0
  
  "00011100","00110010","00101010","00101010","00100110","00011100","00000000","00000000", --1
  "00001000","00001100","00001000","00001000","00001000","00111110","00000000","00000000", --2
  "00011100","00100010","00010000","00001000","00000100","00111110","00000000","00000000", --3
  "00011100","00100010","00010000","00100000","00100010","00011100","00000000","00000000", --4  
  "00011000","00010100","00010010","00111110","00010000","00111100","00000000","00000000", --5
  "00111110","00000010","00111110","00100000","00100010","00011100","00000000","00000000", --6
  "00011100","00100010","00000010","00011110","00100010","00011100","00000000","00000000", --7
  "00111110","00100010","00100000","00010000","00001000","00001000","00000000","00000000", --8
  "00011100","00100010","00011100","00100010","00100010","00011100","00000000","00000000", --9
  "00011100","00100010","00111100","00100000","00100010","00011100","00000000","00000000", --:
  
  "00000000","00001000","00000000","00000000","00000000","00001000","00000000","00000000", --;
  "00000000","00001000","00000000","00000000","00000000","00001000","00001000","00000000", --<
  "00010000","00001000","00000100","00000010","00000100","00001000","00010000","00000000", --=
  "00000000","00000000","00111110","00000000","00000000","00111110","00000000","00000000", -->
  "00000010","00000100","00001000","00010000","00001000","00000100","00000010","00000000", --?
  "00011100","00100010","00011000","00001000","00000000","00001000","00000000","00000000", --@
  "01111100","10000010","10111010","10101010","10111010","10100010","01101100","00000000", --A
  
  "00011100","00100010","00111110","00100010","00100010","00100010","00000000","00000000", --B
  "00011110","00100010","00011110","00100010","00100010","00011110","00000000","00000000", --C
  "00011100","00100010","00000010","00000010","00100010","00011100","00000000","00000000", --D
  "00011110","00100010","00100010","00100010","00100010","00011110","00000000","00000000", --E
  "00111110","00000010","00011110","00000010","00000010","00111110","00000000","00000000", --F
  "00111110","00000010","00011110","00000010","00000010","00000010","00000000","00000000", --G
  "00011100","00100010","00000010","00111010","00100010","00011100","00000000","00000000", --H
  "00100010","00100010","00111110","00100010","00100010","00100010","00000000","00000000", --I
  "00111110","00001000","00001000","00001000","00001000","00111110","00000000","00000000", --J
  "00111000","00010000","00010000","00010000","00010010","00001100","00000000","00000000", --K
  "00010010","00001010","00000110","00001010","00010010","00100010","00000000","00000000", --L
  "00000010","00000010","00000010","00000010","00000010","00111110","00000000","00000000", --M
  "00100010","00110110","00101010","00101010","00100010","00100010","00000000","00000000", --N
  "00100010","00100010","00100110","00101010","00110010","00100010","00000000","00000000", --O
  "00011100","00100010","00100010","00100010","00100010","00011100","00000000","00000000", --P
  "00011110","00100010","00100010","00011110","00000010","00000010","00000000","00000000", --Q
  "00011100","00100010","00100010","00100010","00100010","00011100","01101000","00000000", --R
  "00011110","00100010","00011110","00001010","00010010","00100010","00000000","00000000", --S
  "00111100","00000010","00011100","00100000","00100000","00011110","00000000","00000000", --T
  "00111110","00001000","00001000","00001000","00001000","00001000","00000000","00000000", --U
  "00100010","00100010","00100010","00100010","00100010","00011100","00000000","00000000", --V
  "00100010","00100010","00100010","00010100","00010100","00001000","00000000","00000000", --W
  "00100010","00100010","00100010","00101010","00101010","00010100","00000000","00000000", --X
  "00100010","00010100","00001000","00001000","00010100","00100010","00000000","00000000", --Y
  "00100010","00100010","00011100","00001000","00001000","00001000","00000000","00000000", --Z
  "00111110","00010000","00001000","00000100","00000010","00111110","00000000","00000000", --[
  
  "00011000","00001000","00001000","00001000","00001000","00001000","00011000","00000000", --\
  "00000010","00000100","00001000","00010000","00100000","01000000","00000000","00000000", --]
  "00011000","00010000","00010000","00010000","00010000","00010000","00011000","00000000", --^
  "00001000","00010100","00100010","00000000","00000000","00000000","00000000","00000000", --_
  "00000000","00000000","00000000","00000000","00000000","00000000","11111111","00000000", --`
  "00001000","00010000","00000000","00000000","00000000","00000000","00000000","00000000", --a
  
  "00000000","00011100","00100000","00111100","00100010","01011100","00000000","00000000", --b
  "00000010","00000010","00011010","00100110","00100010","00011110","00000000","00000000", --c
  "00000000","00011100","00000010","00000010","00100010","00011100","00000000","00000000", --d
  "00100000","00100000","00101100","00110010","00100010","00111100","00000000","00000000", --e
  "00000000","00011100","00100010","00111110","00000010","00011100","00000000","00000000", --f
  "00011100","00100010","00000010","00001110","00000010","00000010","00000000","00000000", --g
  "00000000","00111100","00100010","00100010","00111100","00100000","00011100","00000000", --h
  "00000010","00000010","00011010","00100110","00100010","00100010","00000000","00000000", --i
  "00001000","00000000","00001100","00001000","00001000","00011100","00000000","00000000", --j
  "00010000","00000000","00011000","00010000","00010000","00010010","00001100","00000000", --k
  "00000010","00010010","00001010","00001110","00010010","00100010","00000000","00000000", --l
  "00001100","00001000","00001000","00001000","00001000","00111110","00000000","00000000", --m
  "00000000","00010110","00101010","00101010","00101010","00101010","00000000","00000000", --n
  "00000000","00011010","00100100","00100100","00100100","00100100","00000000","00000000", --o
  "00000000","00011100","00100010","00100010","00100010","00011100","00000000","00000000", --p
  "00000000","00011110","00100010","00100010","00011110","00000010","00000010","00000000", --q
  "00000000","00101100","00110010","00100010","00111100","00100000","00100000","00000000", --r
  "00000000","00011010","00100100","00000100","00000100","00000100","00000000","00000000", --s
  "00000000","00111100","00000010","00011100","00100000","00011110","00000000","00000000", --t
  "00000010","00000010","00001110","00000010","00100010","00011100","00000000","00000000", --u
  "00000000","00010010","00010010","00010010","00010010","00101100","00000000","00000000", --v
  "00000000","00100010","00100010","00010100","00010100","00001000","00000000","00000000", --w
  "00000000","00100010","00100010","00101010","00101010","00010100","00000000","00000000", --x
  "00000000","00100010","00010100","00001000","00010100","00100010","00000000","00000000", --y
  "00000000","00100010","00100010","00100010","00111100","00100000","00011100","00000000", --z
  "00000000","00111110","00010000","00001000","00000100","00111110","00000000","00000000", --{
  
  "00010000","00001000","00001000","00000100","00001000","00001000","00010000","00000000", --|
  "00001000","00001000","00001000","00001000","00001000","00001000","00001000","00000000", --}
  "00000100","00001000","00001000","00010000","00001000","00001000","00000100","00000000", --~
  "00000000","00000000","00001100","10010010","01100000","00000000","00000000","00000000", --del
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --0d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --1d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --2d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --3d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --4d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --5d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --6d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --7d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --8d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --9d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --10d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --11d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --12d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --13d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --14d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --15d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --16d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --17d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --18d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --19d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --20d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --21d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --22d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --23d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --24d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --25d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --26d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --27d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --28d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --29d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --30d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --31d
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --space
  
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", --!
  "00001000","00001000","00001000","00001000","00000000","00001000","00000000","00000000", --"
  "00010100","00010100","00000000","00000000","00000000","00000000","00000000","00000000", --#
  "00000000","00010100","00111110","00010100","00111110","00010100","00000000","00000000", --$
  "00001000","00111100","00001010","00011100","00101000","00011110","00001000","00000000", --%
  "10001110","01001010","00101110","00010000","11101000","10100100","11100010","00000000", ----'
  "00001100","00010010","00010010","00001100","00110010","00010010","01101100","00000000", --(
  "00001000","00001000","00000000","00000000","00000000","00000000","00000000","00000000", --)
  "00001000","00000100","00000010","00000010","00000010","00000100","00001000","00000000", --*
  "00001000","00010000","00100000","00100000","00100000","00010000","00001000","00000000", --+
  "00001000","00111110","00010100","00100010","00000000","00000000","00000000","00000000", --,
  "00010000","00010000","00010000","11111110","00010000","00010000","00010000","00000000", ---
  "00000000","00000000","00000000","00000000","00000000","00001000","00001000","00000000", --.
  "00000000","00000000","00000000","00111110","00000000","00000000","00000000","00000000", --/
  "00000000","00000000","00000000","00000000","00000000","00001000","00000000","00000000", --0
  "01000000","00100000","00010000","00001000","00000100","00000010","00000000","00000000", --1
  
  "00011100","00110010","00101010","00101010","00100110","00011100","00000000","00000000", --2
  "00001000","00001100","00001000","00001000","00001000","00111110","00000000","00000000", --3
  "00011100","00100010","00010000","00001000","00000100","00111110","00000000","00000000", --4
  "00011100","00100010","00010000","00100000","00100010","00011100","00000000","00000000", --5
  "00011000","00010100","00010010","00111110","00010000","00111100","00000000","00000000", --6
  "00111110","00000010","00111110","00100000","00100010","00011100","00000000","00000000", --7
  "00011100","00100010","00000010","00011110","00100010","00011100","00000000","00000000", --8
  "00111110","00100010","00100000","00010000","00001000","00001000","00000000","00000000", --9
  "00011100","00100010","00011100","00100010","00100010","00011100","00000000","00000000", --:
  "00011100","00100010","00111100","00100000","00100010","00011100","00000000","00000000", --;
  
  "00000000","00001000","00000000","00000000","00000000","00001000","00000000","00000000", --<
  "00000000","00001000","00000000","00000000","00000000","00001000","00001000","00000000", --=
  "00010000","00001000","00000100","00000010","00000100","00001000","00010000","00000000", -->
  "00000000","00000000","00111110","00000000","00000000","00111110","00000000","00000000", --?
  "00000010","00000100","00001000","00010000","00001000","00000100","00000010","00000000", --@
  "00011100","00100010","00011000","00001000","00000000","00001000","00000000","00000000", --A
  "01111100","10000010","10111010","10101010","10111010","10100010","01101100","00000000", --B
  
  "00011100","00100010","00111110","00100010","00100010","00100010","00000000","00000000", --C
  "00011110","00100010","00011110","00100010","00100010","00011110","00000000","00000000", --D
  "00011100","00100010","00000010","00000010","00100010","00011100","00000000","00000000", --E
  "00011110","00100010","00100010","00100010","00100010","00011110","00000000","00000000", --F
  "00111110","00000010","00011110","00000010","00000010","00111110","00000000","00000000", --G
  "00111110","00000010","00011110","00000010","00000010","00000010","00000000","00000000", --H
  "00011100","00100010","00000010","00111010","00100010","00011100","00000000","00000000", --I
  "00100010","00100010","00111110","00100010","00100010","00100010","00000000","00000000", --J
  "00111110","00001000","00001000","00001000","00001000","00111110","00000000","00000000", --K
  "00111000","00010000","00010000","00010000","00010010","00001100","00000000","00000000", --L
  "00010010","00001010","00000110","00001010","00010010","00100010","00000000","00000000", --M
  "00000010","00000010","00000010","00000010","00000010","00111110","00000000","00000000", --N
  "00100010","00110110","00101010","00101010","00100010","00100010","00000000","00000000", --O
  "00100010","00100010","00100110","00101010","00110010","00100010","00000000","00000000", --P
  "00011100","00100010","00100010","00100010","00100010","00011100","00000000","00000000", --Q
  "00011110","00100010","00100010","00011110","00000010","00000010","00000000","00000000", --R
  "00011100","00100010","00100010","00100010","00100010","00011100","01101000","00000000", --S
  "00011110","00100010","00011110","00001010","00010010","00100010","00000000","00000000", --T
  "00111100","00000010","00011100","00100000","00100000","00011110","00000000","00000000", --U
  "00111110","00001000","00001000","00001000","00001000","00001000","00000000","00000000", --V
  "00100010","00100010","00100010","00100010","00100010","00011100","00000000","00000000", --W
  "00100010","00100010","00100010","00010100","00010100","00001000","00000000","00000000", --X
  "00100010","00100010","00100010","00101010","00101010","00010100","00000000","00000000", --Y
  "00100010","00010100","00001000","00001000","00010100","00100010","00000000","00000000", --Z
  "00100010","00100010","00011100","00001000","00001000","00001000","00000000","00000000", --[
  "00111110","00010000","00001000","00000100","00000010","00111110","00000000","00000000", --\
  
  "00011000","00001000","00001000","00001000","00001000","00001000","00011000","00000000", --]
  "00000010","00000100","00001000","00010000","00100000","01000000","00000000","00000000", --^
  "00011000","00010000","00010000","00010000","00010000","00010000","00011000","00000000", --_
  "00001000","00010100","00100010","00000000","00000000","00000000","00000000","00000000", --`
  "00000000","00000000","00000000","00000000","00000000","00000000","11111111","00000000", --a
  "00001000","00010000","00000000","00000000","00000000","00000000","00000000","00000000", --b
  
  "00000000","00011100","00100000","00111100","00100010","01011100","00000000","00000000", --c
  "00000010","00000010","00011010","00100110","00100010","00011110","00000000","00000000", --d
  "00000000","00011100","00000010","00000010","00100010","00011100","00000000","00000000", --e
  "00100000","00100000","00101100","00110010","00100010","00111100","00000000","00000000", --f
  "00000000","00011100","00100010","00111110","00000010","00011100","00000000","00000000", --g
  "00011100","00100010","00000010","00001110","00000010","00000010","00000000","00000000", --h
  "00000000","00111100","00100010","00100010","00111100","00100000","00011100","00000000", --i
  "00000010","00000010","00011010","00100110","00100010","00100010","00000000","00000000", --j
  "00001000","00000000","00001100","00001000","00001000","00011100","00000000","00000000", --k
  "00010000","00000000","00011000","00010000","00010000","00010010","00001100","00000000", --l
  "00000010","00010010","00001010","00001110","00010010","00100010","00000000","00000000", --m
  "00001100","00001000","00001000","00001000","00001000","00111110","00000000","00000000", --n
  "00000000","00010110","00101010","00101010","00101010","00101010","00000000","00000000", --o
  "00000000","00011010","00100100","00100100","00100100","00100100","00000000","00000000", --p
  "00000000","00011100","00100010","00100010","00100010","00011100","00000000","00000000", --q
  "00000000","00011110","00100010","00100010","00011110","00000010","00000010","00000000", --r
  "00000000","00101100","00110010","00100010","00111100","00100000","00100000","00000000", --s
  "00000000","00011010","00100100","00000100","00000100","00000100","00000000","00000000", --t
  "00000000","00111100","00000010","00011100","00100000","00011110","00000000","00000000", --u
  "00000010","00000010","00001110","00000010","00100010","00011100","00000000","00000000", --v
  "00000000","00010010","00010010","00010010","00010010","00101100","00000000","00000000", --w
  "00000000","00100010","00100010","00010100","00010100","00001000","00000000","00000000", --x
  "00000000","00100010","00100010","00101010","00101010","00010100","00000000","00000000", --y
  "00000000","00100010","00010100","00001000","00010100","00100010","00000000","00000000", --z
  "00000000","00100010","00100010","00100010","00111100","00100000","00011100","00000000", --{
  "00000000","00111110","00010000","00001000","00000100","00111110","00000000","00000000", --|
  
  "00010000","00001000","00001000","00000100","00001000","00001000","00010000","00000000", --}
  "00001000","00001000","00001000","00001000","00001000","00001000","00001000","00000000", --~
  "00000100","00001000","00001000","00010000","00001000","00001000","00000100","00000000", --del
  "00000000","00000000","00001100","10010010","01100000","00000000","00000000","00000000", 
  "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"); 

  component VIDEO_TIME_GEN is
    port ( 
    CLK      : in  Std_logic;
    RST      : in  Std_logic;
    CHARADDR : out Std_logic_vector(12 downto 0);
    PIXROW   : out Std_logic_vector(2 downto 0);
    PIXCOL   : out Std_logic_vector(2 downto 0);
    HSYNCH   : out Std_logic;
    VSYNCH   : out Std_logic;
    BLANK    : out Std_logic);
  end component;

  type CHAR_ARRAY_TYPE is array (0 to 7499)  of Std_logic_vector(7 downto 0);
  signal CHARARRAY : CHAR_ARRAY_TYPE;
  type STATE_TYPE is (GET_COL,ACK_COL,GET_ROW,ACK_ROW,GET_DATA,ACK_DATA);
  signal STATE : STATE_TYPE;

  signal INTHSYNCH, INTVSYNCH   : Std_logic;
  signal HSYNCH_DEL, VSYNCH_DEL : Std_logic;
  signal BLANK, BLANK_DEL, BLANK_DEL_DEL 
                                : Std_logic;
  signal PIX, DATA_WR           : Std_logic;
  signal PIXROW, PIXROW_DEL     : Std_logic_vector(2 downto 0);
  signal PIXCOL, PIXCOL_DEL, PIXCOL_DEL_DEL 
                                : Std_logic_vector(2 downto 0);
  signal CHARADDR               : Std_logic_vector(12 downto 0);
  signal CHAR, PIXELS           : Std_logic_vector(7 downto 0);
  signal ADDRESS                : integer range 0 to 7499;
  signal INT_DATA               : Std_logic_vector(7 downto 0);

begin

  TIMEING1: VIDEO_TIME_GEN port map( 
    CLK      => CLK,
    RST      => RST,
    CHARADDR => CHARADDR, 
    PIXROW   => PIXROW,
    PIXCOL   => PIXCOL,
    HSYNCH   => INTHSYNCH,
    VSYNCH   => INTVSYNCH,
    BLANK    => BLANK
  );

  process
    variable ROW     : integer range 0 to 74;
    variable COL     : integer range 0 to 99;
  begin
    wait until Rising_edge(CLK);
    DATA_WR <= '0';
    case STATE is
      when GET_COL =>
        if DATA_STB = '1' then
          COL := to_integer(unsigned(DATA));
          DATA_ACK <= '1';
          STATE <= ACK_COL;
        end if;
      when ACK_COL =>
        DATA_ACK <= '0';
        STATE <= GET_ROW;
      when GET_ROW =>
        if DATA_STB = '1' then
          ROW := to_integer(unsigned(DATA));
          DATA_ACK <= '1';
          STATE <= ACK_ROW;
        end if;
      when ACK_ROW =>
        DATA_ACK <= '0';
        STATE <= GET_DATA;
      when GET_DATA =>
        if DATA_STB = '1' then
          INT_DATA <= DATA;
          DATA_ACK <= '1';
          STATE <= ACK_DATA;
        end if;
      when ACK_DATA =>
        ADDRESS <= (100*ROW)+COL;
        DATA_WR <= '1';
        DATA_ACK <= '0';
        STATE <= GET_COL;
      when others => null;
    end case;
    if RST = '1' then
      DATA_ACK <= '0';
      STATE <= GET_COL;
    end if;
  end process;

  process(CLK)
  begin
    if Rising_edge(CLK) then
      CHAR <= CHARARRAY(To_integer(Unsigned(CHARADDR)));
      if DATA_WR = '1' then
        CHARARRAY(ADDRESS) <= INT_DATA;
      end if;
    end if; 
  end process;

  process(CLK)
    variable PIXADDRESS :Integer;
    variable PIXVECTOR  : Std_logic_vector(10 downto 0);
  begin
    if Rising_edge(CLK) then
      PIXVECTOR := CHAR & PIXROW_DEL;
      PIXADDRESS := To_integer(Unsigned(PIXVECTOR));
      PIXELS <= PIXARRAY(PIXADDRESS);
    end if;
  end process;

  process(CLK)
  begin
    
    if Rising_edge(CLK) then
      HSYNCH_DEL     <= INTHSYNCH;
      HSYNCH         <= HSYNCH_DEL;
      VSYNCH_DEL     <= INTVSYNCH;
      VSYNCH         <= VSYNCH_DEL;
      BLANK_DEL      <= BLANK;
      BLANK_DEL_DEL  <= BLANK_DEL;
      PIXROW_DEL     <= PIXROW;
      PIXCOL_DEL     <= PIXCOL;
      PIXCOL_DEL_DEL <= PIXCOL_DEL;
    end if;

  end process;

  PIX <= PIXELS(To_integer(Unsigned(PIXCOL_DEL_DEL)));
  
  R <= PIX and not(BLANK_DEL_DEL);
  G <= PIX and not(BLANK_DEL_DEL);
  B <= PIX and not(BLANK_DEL_DEL);
  
end RTL;
  

--+============================================================================+
--|                  *** END OF CHARACTER SVGA DISPLAY ***                     |
--+============================================================================+
