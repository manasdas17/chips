--+============================================================================+
--| +---+----+---+                                              +---+----+---+ |
--| |    \__/    |                                              |    \__/    | |
--|[|            |]--------------------------------------------[|            |]|
--| |            |                                              |            | |
--|[|            |]     This file was generated by Chips       [|            |]|
--| |            |                                              |            | |
--|[|            |]                                            [|            |]|
--| |            |                   Chips                      |            | |
--|[|            |]                                            [|            |]|
--| |            |                                              |            | |
--|[|            |]      http://github.com/dawsonjon/chips     [|            |]|
--| |            |                                              |            | |
--|[|            |]                                            [|            |]|
--| |            |                              Python powered  |            | |
--|[|            |]--------------------------------------------[|            |]|
--| |            |                                              |            | |
--| +------------+                                              +------------+ |
--+============================================================================+

-- generated by python streams library
-- date generated  : UTC 2011-04-20 20:01:33
-- platform        : linux2
-- python version  : 2.6.6 (r266:84292, Sep 15 2010, 16:22:56) [GCC 4.4.5]
-- streams version : 0.1

--+============================================================================+
--|                             **END OF HEADER**                              |
--+============================================================================+

--                                   ***                                       

--+============================================================================+
--|                    **START OF EXTERNAL DEPENDENCIES**                      |
--+============================================================================+


--  ****************************************************************************
--  Filename         :
--  Project          :
--  Version          :0.1
--  Author           :Jonathan P Dawson
--  Created Date     :2005-12-18
--  ****************************************************************************
--  Description      :A RAM based on Xilinx block RAMs
--  ****************************************************************************
--  Dependencies     :Standard Libraries
--  ****************************************************************************
--  Revision History :
--  
--  Date :2005-12-18
--  Author :Jonathan P Dawson
--  Modification: Created File
--  
--  ****************************************************************************
--  Copyright (C) Jonathan P Dawson 2005
--  ****************************************************************************
 library ieee;
 use ieee.std_logic_1164.all;
 use ieee.numeric_std.all;

 entity RAMARRAY is
    generic(
        DEPTH : integer;
        WIDTH : integer
    );
    port(
        CLK             : in  std_logic;
        RST             : in  std_logic;
        ADDRESS_IN      : in  std_logic_vector;
        ADDRESS_IN_STB  : in  std_logic;
        ADDRESS_IN_ACK  : out std_logic;
        DATA_IN         : in  std_logic_vector;
        DATA_IN_STB     : in  std_logic;
        DATA_IN_ACK     : out std_logic;
        ADDRESS_OUT     : in  std_logic_vector;
        ADDRESS_OUT_STB : in  std_logic;
        ADDRESS_OUT_ACK : out std_logic;
        DATA_OUT        : out std_logic_vector;
        DATA_OUT_STB    : out std_logic;
        DATA_OUT_ACK    : in  std_logic
    );
  end entity RAMARRAY;

  architecture RTL of RAMARRAY is

    type MEMORY_TYPE is array (0 to DEPTH-1) of std_logic_vector(WIDTH-1 downto 0);
    shared variable MEMORY : MEMORY_TYPE;

    type IN_STATE_TYPE is (READ_IN_ADDRESS, ACK_IN_ADDRESS, READ_IN_DATA, ACK_IN_DATA);
    signal IN_STATE : IN_STATE_TYPE;

    type OUT_STATE_TYPE is (READ_OUT_ADDRESS, ACK_OUT_ADDRESS, WRITE_OUT_DATA);
    signal OUT_STATE : OUT_STATE_TYPE;

  begin

     process
      variable ADDRESS : integer range 0 to DEPTH-1;
    begin
      wait until rising_edge(CLK);
      case IN_STATE is

        when READ_IN_ADDRESS =>
           if ADDRESS_IN_STB = '1' then
               ADDRESS := to_integer(unsigned(ADDRESS_IN));
               ADDRESS_IN_ACK <= '1';
               IN_STATE <= ACK_IN_ADDRESS;
           end if;

        when ACK_IN_ADDRESS =>
           ADDRESS_IN_ACK <= '0';
           IN_STATE <= READ_IN_DATA;

        when READ_IN_DATA =>
           if DATA_IN_STB = '1' then
               MEMORY(ADDRESS) := DATA_IN;
               DATA_IN_ACK <= '1';
               IN_STATE <= ACK_IN_DATA;
           end if;

        when ACK_IN_DATA =>
           DATA_IN_ACK <= '0';
           IN_STATE <= READ_IN_ADDRESS;

        when others => IN_STATE <= READ_IN_ADDRESS;

      end case;
      if RST = '1' then
        DATA_IN_ACK <= '0';
        ADDRESS_IN_ACK <= '0';
        IN_STATE <= READ_IN_ADDRESS;
      end if;
    end process;

    process
       variable ADDRESS : integer range 0 to DEPTH-1;
    begin
      wait until rising_edge(CLK);
      case OUT_STATE is

        when READ_OUT_ADDRESS =>
           if ADDRESS_OUT_STB = '1' then
             ADDRESS := to_integer(unsigned(ADDRESS_OUT));
             ADDRESS_OUT_ACK <= '1';
             OUT_STATE <= ACK_OUT_ADDRESS;
           end if;

        when ACK_OUT_ADDRESS =>
           ADDRESS_OUT_ACK <= '0';
           OUT_STATE <= WRITE_OUT_DATA;

        when WRITE_OUT_DATA =>
           DATA_OUT <= MEMORY(ADDRESS);
           DATA_OUT_STB <= '1';
           if DATA_OUT_ACK = '1' then
             DATA_OUT_STB <= '0';
             OUT_STATE <= READ_OUT_ADDRESS;
           end if;

        when others => OUT_STATE <= READ_OUT_ADDRESS;

      end case;
      if RST = '1' then
        DATA_OUT_STB <= '0';
        ADDRESS_OUT_ACK <= '0';
        OUT_STATE <= READ_OUT_ADDRESS;
      end if;
  end process;

end RTL;
--  ****************************************************************************
--  End of RAM
--  ****************************************************************************

--+============================================================================+
--|                     **END OF EXTERNAL DEPENDENCIES**                       |
--+============================================================================+

--                                   ***                                       

--+============================================================================+
--|                     **START OF AUTO GENERATED CODE**                       |
--+============================================================================+

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity STREAMS_VHDL_MODEL is

end entity STREAMS_VHDL_MODEL;

architecture RTL of STREAMS_VHDL_MODEL is


  --returns the greater of the two parameters
  function MAX(
    A : integer;
    B : integer) return integer is
  begin
    if A > B then
      return A;
    else
      return B;
    end if;
  end MAX;

  --returns a std_logic_vector sum of the two parameters
  function ABSOLUTE(
    A : std_logic_vector) return std_logic_vector is
  begin
    return std_logic_vector(abs(signed(A)));
  end ABSOLUTE;

  --returns a std_logic_vector sum of the two parameters
  function ADD(
    A : std_logic_vector; 
    B : std_logic_vector) return std_logic_vector is
  begin
    return std_logic_vector(
      resize(signed(A), MAX(A'length, B'length) + 1) + 
      resize(signed(B), MAX(A'length, B'length) + 1));
    end ADD;

  --returns a std_logic_vector product of the two parameters
  function MUL(
    A : std_logic_vector; 
    B : std_logic_vector) return std_logic_vector is
  begin
    return std_logic_vector(
      signed(A) *
      signed(B));
    end MUL;

  --returns a std_logic_vector difference of the two parameters
  function SUB(
    A : std_logic_vector; 
    B : std_logic_vector) return std_logic_vector is
  begin
    return std_logic_vector(
      resize(signed(A), MAX(A'length, B'length) + 1) - 
      resize(signed(B), MAX(A'length, B'length) + 1));
  end SUB;

  --returns A shifted right (arithmetic) by A
  function SR(
    A  : std_logic_vector; 
    B : std_logic_vector) return std_logic_vector is
  begin
    return std_logic_vector(shift_right(signed(A), to_integer(signed(B))));
  end SR;

  --returns A shifted left by B
  function SL(
    A  : std_logic_vector; 
    B : std_logic_vector) return std_logic_vector is
  begin
    return std_logic_vector(shift_left(signed(A), to_integer(signed(B))));
  end SL;

  --returns bitwise and of A and B
  --(A and B are resized to the length of the larger first)
  function BAND(
    A : std_logic_vector; 
    B : std_logic_vector) return std_logic_vector is
  begin
    return std_logic_vector(
      resize(signed(A), MAX(A'LENGTH, B'LENGTH)) and
      resize(signed(B), MAX(A'LENGTH, B'LENGTH)));
  end BAND;

  --returns bitwise or of A and B
  --(A and B are resized to the length of the larger first)
  function BOR(
    A : std_logic_vector; 
    B : std_logic_vector) return std_logic_vector is
  begin
    return std_logic_vector(
      resize(signed(A), MAX(A'LENGTH, B'LENGTH)) or
      resize(signed(B), MAX(A'LENGTH, B'LENGTH)));
  end BOR;

  --returns bitwise xor of A and B
  --(A and B are resized to the length of the larger first)
  function BXOR(
    A : std_logic_vector; 
    B : std_logic_vector) return std_logic_vector is
  begin
    return std_logic_vector(
      resize(signed(A), MAX(A'LENGTH, B'LENGTH)) xor
      resize(signed(B), MAX(A'LENGTH, B'LENGTH)));
  end BXOR;

  --equality comparison of A and B
  --(A and B are resized to the length of the larger first)
  function EQ(
    A : std_logic_vector; 
    B : std_logic_vector) return std_logic_vector is
  begin
    if 
      resize(signed(A), MAX(A'LENGTH, B'LENGTH)) =
      resize(signed(B), MAX(A'LENGTH, B'LENGTH)) then
      return "1";
    else
      return "0";
    end if;
  end EQ;

  --inequality comparison of A and B
  --(A and B are resized to the length of the larger first)
  function NE(
    A : std_logic_vector; 
    B : std_logic_vector) return std_logic_vector is
  begin
    if 
    resize(signed(A), MAX(A'LENGTH, B'LENGTH)) /=
    resize(signed(B), MAX(A'LENGTH, B'LENGTH)) then
      return "1";
    else
      return "0";
    end if;
  end NE;

  --greater than comparison of A and B
  --(A and B are resized to the length of the larger first)
  function GT(
    A : std_logic_vector; 
    B : std_logic_vector) return std_logic_vector is
  begin
    if 
      resize(signed(A), MAX(A'LENGTH, B'LENGTH)) >
      resize(signed(B), MAX(A'LENGTH, B'LENGTH)) then
      return "1";
    else
      return "0";
    end if;
  end GT;

  --greater than or equal comparison of A and B
  --(A and B are resized to the length of the larger first)
  function GE(
    A : std_logic_vector; 
    B : std_logic_vector) return std_logic_vector is
  begin
    if 
      resize(signed(A), MAX(A'LENGTH, B'LENGTH)) >=
      resize(signed(B), MAX(A'LENGTH, B'LENGTH)) then
      return "1";
    else
      return "0";
    end if;
  end GE;

  --less than comparison of A and B
  --(A and B are resized to the length of the larger first)
  function LT(
    A : std_logic_vector; 
    B : std_logic_vector) return std_logic_vector is
  begin
    if 
      resize(signed(A), MAX(A'LENGTH, B'LENGTH)) <
      resize(signed(B), MAX(A'LENGTH, B'LENGTH)) then
      return "1";
    else
      return "0";
    end if;
  end LT;

  --less than or equal comparison of A and B
  --(A and B are resized to the length of the larger first)
  function LE(
    A : std_logic_vector; 
    B : std_logic_vector) return std_logic_vector is
  begin
    if 
      resize(signed(A), MAX(A'LENGTH, B'LENGTH)) <=
      resize(signed(B), MAX(A'LENGTH, B'LENGTH)) then
      return "1";
    else
      return "0";
    end if;
  end LE;

  --logical negation
  function LNOT(
    A : std_logic_vector) return std_logic_vector is
  begin
    if 
      A = std_logic_vector(to_signed(0, A'LENGTH)) then
      return "1";
    else
      return "0";
    end if;
  end LNOT;

  --resize A to B bits
  function STD_RESIZE(
    A : std_logic_vector; 
    B : integer) return std_logic_vector is
  begin
    return std_logic_vector(
      resize(signed(A), B));
  end STD_RESIZE;

  type BINARY_STATE_TYPE is (BINARY_INPUT, BINARY_OUTPUT);
  type UNARY_STATE_TYPE is (UNARY_INPUT, UNARY_OUTPUT);
  type TEE_STATE_TYPE is (TEE_INPUT_A, TEE_WAIT_YZ, TEE_WAIT_Y, TEE_WAIT_Z);
  type DIVIDER_STATE_TYPE is (READ_A_B, DIVIDE_1, DIVIDE_2, WRITE_Z);
  type SERIAL_IN_STATE_TYPE is (IDLE, START, RX0, RX1, RX2, RX3, RX4, RX5, RX6, RX7, STOP, OUTPUT_DATA);
  type SERIAL_OUT_STATE_TYPE is (IDLE, START, WAIT_EN, TX0, TX1, TX2, TX3, TX4, TX5, TX6, TX7, STOP);
  type PRINTER_STATE_TYPE is (INPUT_A, SHIFT, OUTPUT_SIGN, OUTPUT_Z, OUTPUT_NL);
  type HEX_PRINTER_STATE_TYPE is (INPUT_A, OUTPUT_SIGN, OUTPUT_DIGITS);

  constant TIMER_1us_MAX : integer := 49;
  signal TIMER_1us_COUNT : integer range 0 to TIMER_1us_MAX;
  signal TIMER_1us : std_logic;
  constant TIMER_10us_MAX : integer := 49;
  signal TIMER_10us_COUNT : integer range 0 to TIMER_1us_MAX;
  signal TIMER_10us : std_logic;
  constant TIMER_100us_MAX : integer := 49;
  signal TIMER_100us_COUNT : integer range 0 to TIMER_1us_MAX;
  signal TIMER_100us : std_logic;
  constant TIMER_1ms_MAX : integer := 49;
  signal TIMER_1ms_COUNT : integer range 0 to TIMER_1us_MAX;
  signal TIMER_1ms : std_logic;

  signal CLK : std_logic;
  signal RST : std_logic;
  signal STREAM_1     : std_logic_vector(8 downto 0);
  signal STREAM_1_STB : std_logic;
  signal STREAM_1_ACK : std_logic;
  signal STATE_1 : UNARY_STATE_TYPE;
  type LOOKUP_1_TYPE is array (0 to 16383) of std_logic_vector(8 downto 0);
  signal LOOKUP_1 : LOOKUP_1_TYPE := (
0 => "001100110",
1 => "001100110",
2 => "001100111",
3 => "001100101",
4 => "001100111",
5 => "001101000",
6 => "001101001",
7 => "001101000",
8 => "001101000",
9 => "001101011",
10 => "001101011",
11 => "001101100",
12 => "001101100",
13 => "001101101",
14 => "001101110",
15 => "001101111",
16 => "001110000",
17 => "001101111",
18 => "001101110",
19 => "001101100",
20 => "001101011",
21 => "001101100",
22 => "001101011",
23 => "001101100",
24 => "001101101",
25 => "001101101",
26 => "001101101",
27 => "001101111",
28 => "001101111",
29 => "001110001",
30 => "001101110",
31 => "001101111",
32 => "001101111",
33 => "001101111",
34 => "001101101",
35 => "001101110",
36 => "001101110",
37 => "001101100",
38 => "001101110",
39 => "001101100",
40 => "001101101",
41 => "001101101",
42 => "001101010",
43 => "001101010",
44 => "001101110",
45 => "001101111",
46 => "001101111",
47 => "001101100",
48 => "001101111",
49 => "001101110",
50 => "001110000",
51 => "001101101",
52 => "001101110",
53 => "001101101",
54 => "001101001",
55 => "001101100",
56 => "001101010",
57 => "001101100",
58 => "001101011",
59 => "001101011",
60 => "001101101",
61 => "001101011",
62 => "001101101",
63 => "001101111",
64 => "001101101",
65 => "001101100",
66 => "001101011",
67 => "001101011",
68 => "001101011",
69 => "001101001",
70 => "001101010",
71 => "001101011",
72 => "001101010",
73 => "001100111",
74 => "001101100",
75 => "001101100",
76 => "001101110",
77 => "001101101",
78 => "001101101",
79 => "001101011",
80 => "001101101",
81 => "001101011",
82 => "001101001",
83 => "001100110",
84 => "001100100",
85 => "001100011",
86 => "001100101",
87 => "001100111",
88 => "001101000",
89 => "001100101",
90 => "001101000",
91 => "001101000",
92 => "001100110",
93 => "001100101",
94 => "001100001",
95 => "001100010",
96 => "001100100",
97 => "001100101",
98 => "001100011",
99 => "001100000",
100 => "001100010",
101 => "001100100",
102 => "001100100",
103 => "001100101",
104 => "001100000",
105 => "001100001",
106 => "001100001",
107 => "001100001",
108 => "001100100",
109 => "001100010",
110 => "001100100",
111 => "001100100",
112 => "001100000",
113 => "001100101",
114 => "001011111",
115 => "001011111",
116 => "001100001",
117 => "001011110",
118 => "001011111",
119 => "001011101",
120 => "001011110",
121 => "001011110",
122 => "001011110",
123 => "001011100",
124 => "001011011",
125 => "001011011",
126 => "001010111",
127 => "001011100",
128 => "001100101",
129 => "001101000",
130 => "001101000",
131 => "001101100",
132 => "001101010",
133 => "001101011",
134 => "001101000",
135 => "001101000",
136 => "001101000",
137 => "001101000",
138 => "001101011",
139 => "001101011",
140 => "001101100",
141 => "001101011",
142 => "001101011",
143 => "001101011",
144 => "001101011",
145 => "001101001",
146 => "001101011",
147 => "001101010",
148 => "001101001",
149 => "001101000",
150 => "001101010",
151 => "001101010",
152 => "001101010",
153 => "001101010",
154 => "001101001",
155 => "001101011",
156 => "001101011",
157 => "001101010",
158 => "001101101",
159 => "001101111",
160 => "001101011",
161 => "001101101",
162 => "001101101",
163 => "001101111",
164 => "001101101",
165 => "001101111",
166 => "001101100",
167 => "001101100",
168 => "001110000",
169 => "001110001",
170 => "001110001",
171 => "001110001",
172 => "001110001",
173 => "001101111",
174 => "001110001",
175 => "001101110",
176 => "001101111",
177 => "001101110",
178 => "001101101",
179 => "001101110",
180 => "001101110",
181 => "001101101",
182 => "001101100",
183 => "001101100",
184 => "001101100",
185 => "001101111",
186 => "001101010",
187 => "001101011",
188 => "001101010",
189 => "001101010",
190 => "001101010",
191 => "001101011",
192 => "001101101",
193 => "001101100",
194 => "001101110",
195 => "001101111",
196 => "001101101",
197 => "001101001",
198 => "001101000",
199 => "001101100",
200 => "001101111",
201 => "001101101",
202 => "001101101",
203 => "001101110",
204 => "001101110",
205 => "001101101",
206 => "001101011",
207 => "001101000",
208 => "001101000",
209 => "001101001",
210 => "001101000",
211 => "001100010",
212 => "001100010",
213 => "001100101",
214 => "001100101",
215 => "001100110",
216 => "001101010",
217 => "001101011",
218 => "001101011",
219 => "001101100",
220 => "001101000",
221 => "001100101",
222 => "001100110",
223 => "001100101",
224 => "001011111",
225 => "001100011",
226 => "001100100",
227 => "001100110",
228 => "001100111",
229 => "001100110",
230 => "001100010",
231 => "001100011",
232 => "001100000",
233 => "001100001",
234 => "001100010",
235 => "001100001",
236 => "001100001",
237 => "001100010",
238 => "001100010",
239 => "001100010",
240 => "001100001",
241 => "001011110",
242 => "001011111",
243 => "001100000",
244 => "001100001",
245 => "001100000",
246 => "001011100",
247 => "001011011",
248 => "001011100",
249 => "001011010",
250 => "001011110",
251 => "001011001",
252 => "001011110",
253 => "001011110",
254 => "001011010",
255 => "001011011",
256 => "001101001",
257 => "001101101",
258 => "001101100",
259 => "001101100",
260 => "001101010",
261 => "001101011",
262 => "001101011",
263 => "001101101",
264 => "001101010",
265 => "001101001",
266 => "001101011",
267 => "001101011",
268 => "001101000",
269 => "001101011",
270 => "001101010",
271 => "001101010",
272 => "001101001",
273 => "001101010",
274 => "001100110",
275 => "001100100",
276 => "001101100",
277 => "001101111",
278 => "001101110",
279 => "001101100",
280 => "001101011",
281 => "001101110",
282 => "001101110",
283 => "001110000",
284 => "001110000",
285 => "001101101",
286 => "001101101",
287 => "001101110",
288 => "001101100",
289 => "001101101",
290 => "001101100",
291 => "001101011",
292 => "001101100",
293 => "001101101",
294 => "001101011",
295 => "001101100",
296 => "001101011",
297 => "001101101",
298 => "001101011",
299 => "001101110",
300 => "001101101",
301 => "001101101",
302 => "001101001",
303 => "001101001",
304 => "001101000",
305 => "001101110",
306 => "001101100",
307 => "001101011",
308 => "001101000",
309 => "001101110",
310 => "001101101",
311 => "001101110",
312 => "001110001",
313 => "001101011",
314 => "001101011",
315 => "001101111",
316 => "001101101",
317 => "001101100",
318 => "001101101",
319 => "001110000",
320 => "001101101",
321 => "001110000",
322 => "001101110",
323 => "001101011",
324 => "001101101",
325 => "001101011",
326 => "001101001",
327 => "001101100",
328 => "001101011",
329 => "001101101",
330 => "001101010",
331 => "001101011",
332 => "001101011",
333 => "001101001",
334 => "001100111",
335 => "001101001",
336 => "001101011",
337 => "001101100",
338 => "001101010",
339 => "001101011",
340 => "001101001",
341 => "001100101",
342 => "001101001",
343 => "001100101",
344 => "001100111",
345 => "001101100",
346 => "001101010",
347 => "001101001",
348 => "001101001",
349 => "001101000",
350 => "001101001",
351 => "001100110",
352 => "001100101",
353 => "001100110",
354 => "001100101",
355 => "001100011",
356 => "001100101",
357 => "001100010",
358 => "001100111",
359 => "001100101",
360 => "001100010",
361 => "001100001",
362 => "001100001",
363 => "001100000",
364 => "001011110",
365 => "001100010",
366 => "001100000",
367 => "001011100",
368 => "001011110",
369 => "001011101",
370 => "001011111",
371 => "001100001",
372 => "001011111",
373 => "001011100",
374 => "001011000",
375 => "001011011",
376 => "001011100",
377 => "001011100",
378 => "001011100",
379 => "001011000",
380 => "001011010",
381 => "001011010",
382 => "001011110",
383 => "001011110",
384 => "001100101",
385 => "001100110",
386 => "001101000",
387 => "001101011",
388 => "001101011",
389 => "001101101",
390 => "001101101",
391 => "001101010",
392 => "001100111",
393 => "001100100",
394 => "001101001",
395 => "001101001",
396 => "001101001",
397 => "001101010",
398 => "001101011",
399 => "001101000",
400 => "001101100",
401 => "001101010",
402 => "001101011",
403 => "001101100",
404 => "001101100",
405 => "001101110",
406 => "001101110",
407 => "001101111",
408 => "001101110",
409 => "001101111",
410 => "001101110",
411 => "001101110",
412 => "001110001",
413 => "001101111",
414 => "001101100",
415 => "001101011",
416 => "001101110",
417 => "001101110",
418 => "001101100",
419 => "001101011",
420 => "001101101",
421 => "001101011",
422 => "001101110",
423 => "001101100",
424 => "001101101",
425 => "001101111",
426 => "001101100",
427 => "001101110",
428 => "001110001",
429 => "001110000",
430 => "001101110",
431 => "001101101",
432 => "001101111",
433 => "001101111",
434 => "001101100",
435 => "001101101",
436 => "001101110",
437 => "001101101",
438 => "001101101",
439 => "001110000",
440 => "001101101",
441 => "001101110",
442 => "001101011",
443 => "001101110",
444 => "001101111",
445 => "001101010",
446 => "001101101",
447 => "001101011",
448 => "001100111",
449 => "001101000",
450 => "001101001",
451 => "001101010",
452 => "001101010",
453 => "001101010",
454 => "001101010",
455 => "001100111",
456 => "001100110",
457 => "001101100",
458 => "001101110",
459 => "001101101",
460 => "001101010",
461 => "001101011",
462 => "001100110",
463 => "001100110",
464 => "001100100",
465 => "001101101",
466 => "001101011",
467 => "001101111",
468 => "001101100",
469 => "001101011",
470 => "001101001",
471 => "001101010",
472 => "001101000",
473 => "001100100",
474 => "001100010",
475 => "001100100",
476 => "001100101",
477 => "001101000",
478 => "001100110",
479 => "001101010",
480 => "001100101",
481 => "001100011",
482 => "001100101",
483 => "001100101",
484 => "001101000",
485 => "001100110",
486 => "001100111",
487 => "001100110",
488 => "001100101",
489 => "001100101",
490 => "001100010",
491 => "001011111",
492 => "001100000",
493 => "001100000",
494 => "001100000",
495 => "001100010",
496 => "001011101",
497 => "001011111",
498 => "001011110",
499 => "001011111",
500 => "001011010",
501 => "001011010",
502 => "001011100",
503 => "001011001",
504 => "001011010",
505 => "001011111",
506 => "001100000",
507 => "001011101",
508 => "001011100",
509 => "001100100",
510 => "001100011",
511 => "001100110",
512 => "001100101",
513 => "001100101",
514 => "001100101",
515 => "001100101",
516 => "001101001",
517 => "001101001",
518 => "001101010",
519 => "001101010",
520 => "001101100",
521 => "001101110",
522 => "001101001",
523 => "001100100",
524 => "001101010",
525 => "001101000",
526 => "001100110",
527 => "001100111",
528 => "001101001",
529 => "001101001",
530 => "001101011",
531 => "001101011",
532 => "001101101",
533 => "001101100",
534 => "001101011",
535 => "001101011",
536 => "001101110",
537 => "001101101",
538 => "001101110",
539 => "001101100",
540 => "001101011",
541 => "001101101",
542 => "001101000",
543 => "001101101",
544 => "001101100",
545 => "001101110",
546 => "001101100",
547 => "001101111",
548 => "001101110",
549 => "001101101",
550 => "001101110",
551 => "001101110",
552 => "001110000",
553 => "001101111",
554 => "001101101",
555 => "001101110",
556 => "001101101",
557 => "001110001",
558 => "001110010",
559 => "001101110",
560 => "001101111",
561 => "001101110",
562 => "001101110",
563 => "001101100",
564 => "001110010",
565 => "001101110",
566 => "001110000",
567 => "001101110",
568 => "001101110",
569 => "001101010",
570 => "001101011",
571 => "001101000",
572 => "001101001",
573 => "001101001",
574 => "001101000",
575 => "001101001",
576 => "001100110",
577 => "001101001",
578 => "001100101",
579 => "001100111",
580 => "001100101",
581 => "001100100",
582 => "001100101",
583 => "001100110",
584 => "001100101",
585 => "001100111",
586 => "001101010",
587 => "001101001",
588 => "001101100",
589 => "001101010",
590 => "001101011",
591 => "001101101",
592 => "001101001",
593 => "001101011",
594 => "001101001",
595 => "001101011",
596 => "001101010",
597 => "001101010",
598 => "001101100",
599 => "001101001",
600 => "001101001",
601 => "001101000",
602 => "001101000",
603 => "001100010",
604 => "001101000",
605 => "001101001",
606 => "001100100",
607 => "001011111",
608 => "001100101",
609 => "001100100",
610 => "001100011",
611 => "001100110",
612 => "001100110",
613 => "001100111",
614 => "001100111",
615 => "001100110",
616 => "001100100",
617 => "001100110",
618 => "001100100",
619 => "001100000",
620 => "001100011",
621 => "001100011",
622 => "001100000",
623 => "001011110",
624 => "001100100",
625 => "001100001",
626 => "001011100",
627 => "001011111",
628 => "001011110",
629 => "001011111",
630 => "001011110",
631 => "001100000",
632 => "001011101",
633 => "001100001",
634 => "001100010",
635 => "001011101",
636 => "001100011",
637 => "001100101",
638 => "001101110",
639 => "001101111",
640 => "001100011",
641 => "001100101",
642 => "001100101",
643 => "001100011",
644 => "001100010",
645 => "001101001",
646 => "001101000",
647 => "001101000",
648 => "001101001",
649 => "001101010",
650 => "001101100",
651 => "001101011",
652 => "001101010",
653 => "001101010",
654 => "001101001",
655 => "001101011",
656 => "001101010",
657 => "001101000",
658 => "001100111",
659 => "001101100",
660 => "001101101",
661 => "001101001",
662 => "001101100",
663 => "001101010",
664 => "001101100",
665 => "001101100",
666 => "001101101",
667 => "001101011",
668 => "001101101",
669 => "001101101",
670 => "001101100",
671 => "001101100",
672 => "001101011",
673 => "001101110",
674 => "001101110",
675 => "001101111",
676 => "001101101",
677 => "001101101",
678 => "001101111",
679 => "001110000",
680 => "001110001",
681 => "001110001",
682 => "001101110",
683 => "001101111",
684 => "001101101",
685 => "001101111",
686 => "001101101",
687 => "001101110",
688 => "001101101",
689 => "001110000",
690 => "001101101",
691 => "001101111",
692 => "001101011",
693 => "001101010",
694 => "001101001",
695 => "001101011",
696 => "001101011",
697 => "001101001",
698 => "001101010",
699 => "001101010",
700 => "001100110",
701 => "001101001",
702 => "001101011",
703 => "001101011",
704 => "001101000",
705 => "001100100",
706 => "001100111",
707 => "001100111",
708 => "001100101",
709 => "001100100",
710 => "001100100",
711 => "001100101",
712 => "001101000",
713 => "001101001",
714 => "001100110",
715 => "001101010",
716 => "001101001",
717 => "001101101",
718 => "001101001",
719 => "001101101",
720 => "001101111",
721 => "001110001",
722 => "001110000",
723 => "001101110",
724 => "001110000",
725 => "001101110",
726 => "001101010",
727 => "001101100",
728 => "001101100",
729 => "001101001",
730 => "001101010",
731 => "001101001",
732 => "001101101",
733 => "001101011",
734 => "001100111",
735 => "001101001",
736 => "001100000",
737 => "001011111",
738 => "001100001",
739 => "001011111",
740 => "001011011",
741 => "001100001",
742 => "001100010",
743 => "001100100",
744 => "001100101",
745 => "001100000",
746 => "001100011",
747 => "001011111",
748 => "001011100",
749 => "001011010",
750 => "001100000",
751 => "001100000",
752 => "001100100",
753 => "001100010",
754 => "001100011",
755 => "001100010",
756 => "001100101",
757 => "001100101",
758 => "001100111",
759 => "001100111",
760 => "001101010",
761 => "001101000",
762 => "001101001",
763 => "001101100",
764 => "001110000",
765 => "001110001",
766 => "001110101",
767 => "001101111",
768 => "001100010",
769 => "001100010",
770 => "001100101",
771 => "001100101",
772 => "001101000",
773 => "001100111",
774 => "001101001",
775 => "001101000",
776 => "001101010",
777 => "001101100",
778 => "001101100",
779 => "001101010",
780 => "001101011",
781 => "001101001",
782 => "001100011",
783 => "001100100",
784 => "001101001",
785 => "001100111",
786 => "001101010",
787 => "001101011",
788 => "001101001",
789 => "001101001",
790 => "001101000",
791 => "001100111",
792 => "001100100",
793 => "001100100",
794 => "001100110",
795 => "001101010",
796 => "001101100",
797 => "001101110",
798 => "001101000",
799 => "001101001",
800 => "001101100",
801 => "001101001",
802 => "001101010",
803 => "001101101",
804 => "001101110",
805 => "001101110",
806 => "001110000",
807 => "001101110",
808 => "001101100",
809 => "001101110",
810 => "001101011",
811 => "001101010",
812 => "001101100",
813 => "001101101",
814 => "001101000",
815 => "001101011",
816 => "001101011",
817 => "001101010",
818 => "001101110",
819 => "001101010",
820 => "001101011",
821 => "001101001",
822 => "001100111",
823 => "001101100",
824 => "001101000",
825 => "001101011",
826 => "001101100",
827 => "001101010",
828 => "001101011",
829 => "001101000",
830 => "001101001",
831 => "001101010",
832 => "001100111",
833 => "001100111",
834 => "001100111",
835 => "001100111",
836 => "001101000",
837 => "001100110",
838 => "001100111",
839 => "001100101",
840 => "001011110",
841 => "001100100",
842 => "001100110",
843 => "001011111",
844 => "001100111",
845 => "001101011",
846 => "001100110",
847 => "001100111",
848 => "001101000",
849 => "001100110",
850 => "001101001",
851 => "001100111",
852 => "001101110",
853 => "001101110",
854 => "001101100",
855 => "001101011",
856 => "001100101",
857 => "001100110",
858 => "001100100",
859 => "001100010",
860 => "001101010",
861 => "001101011",
862 => "001100111",
863 => "001100000",
864 => "001011111",
865 => "001011101",
866 => "001011111",
867 => "001011111",
868 => "001100010",
869 => "001100011",
870 => "001100010",
871 => "001100100",
872 => "001100010",
873 => "001100001",
874 => "001100000",
875 => "001100011",
876 => "001100011",
877 => "001101001",
878 => "001101010",
879 => "001100110",
880 => "001100111",
881 => "001110100",
882 => "001101011",
883 => "001100010",
884 => "001100001",
885 => "001110011",
886 => "001110000",
887 => "001110000",
888 => "001110111",
889 => "001110010",
890 => "001101111",
891 => "001110011",
892 => "001110000",
893 => "001101001",
894 => "001101000",
895 => "001101001",
896 => "001011111",
897 => "001100001",
898 => "001011111",
899 => "001100000",
900 => "001100000",
901 => "001100101",
902 => "001100110",
903 => "001101000",
904 => "001100111",
905 => "001101011",
906 => "001101110",
907 => "001101100",
908 => "001101100",
909 => "001101010",
910 => "001100111",
911 => "001101001",
912 => "001101011",
913 => "001101001",
914 => "001101001",
915 => "001101100",
916 => "001101010",
917 => "001101011",
918 => "001101101",
919 => "001101100",
920 => "001101011",
921 => "001101000",
922 => "001100011",
923 => "001101010",
924 => "001101001",
925 => "001101101",
926 => "001101101",
927 => "001101111",
928 => "001101101",
929 => "001101010",
930 => "001100100",
931 => "001101100",
932 => "001101110",
933 => "001101110",
934 => "001101111",
935 => "001101010",
936 => "001101011",
937 => "001101101",
938 => "001101001",
939 => "001100110",
940 => "001100101",
941 => "001101010",
942 => "001100101",
943 => "001100110",
944 => "001100110",
945 => "001100110",
946 => "001101010",
947 => "001101010",
948 => "001101010",
949 => "001101110",
950 => "001101110",
951 => "001101110",
952 => "001101100",
953 => "001110000",
954 => "001110000",
955 => "001110000",
956 => "001101100",
957 => "001101111",
958 => "001110011",
959 => "001110000",
960 => "001101111",
961 => "001101101",
962 => "001101100",
963 => "001101100",
964 => "001101100",
965 => "001101010",
966 => "001101001",
967 => "001100111",
968 => "001101011",
969 => "001101001",
970 => "001100110",
971 => "001101011",
972 => "001101000",
973 => "001100111",
974 => "001101000",
975 => "001100110",
976 => "001100111",
977 => "001101101",
978 => "001101101",
979 => "001101010",
980 => "001100110",
981 => "001101000",
982 => "001101001",
983 => "001100110",
984 => "001100110",
985 => "001100101",
986 => "001100010",
987 => "001101100",
988 => "001101000",
989 => "001101001",
990 => "001100100",
991 => "001101001",
992 => "001100111",
993 => "001100100",
994 => "001100101",
995 => "001100110",
996 => "001100101",
997 => "001100010",
998 => "001101000",
999 => "001100111",
1000 => "001101101",
1001 => "001101101",
1002 => "001110111",
1003 => "001110100",
1004 => "001101111",
1005 => "001110101",
1006 => "001110010",
1007 => "001110000",
1008 => "001101101",
1009 => "001101111",
1010 => "001100111",
1011 => "001100110",
1012 => "001100010",
1013 => "001101010",
1014 => "001110000",
1015 => "001101011",
1016 => "001101101",
1017 => "001101111",
1018 => "001110000",
1019 => "001100110",
1020 => "001101000",
1021 => "001101001",
1022 => "001100100",
1023 => "001100010",
1024 => "001100100",
1025 => "001100000",
1026 => "001100001",
1027 => "001100100",
1028 => "001100000",
1029 => "001100110",
1030 => "001101001",
1031 => "001101010",
1032 => "001101000",
1033 => "001100111",
1034 => "001101010",
1035 => "001100111",
1036 => "001101001",
1037 => "001101001",
1038 => "001101001",
1039 => "001101010",
1040 => "001101010",
1041 => "001101001",
1042 => "001101100",
1043 => "001100110",
1044 => "001101000",
1045 => "001101011",
1046 => "001101100",
1047 => "001101111",
1048 => "001101100",
1049 => "001101100",
1050 => "001101001",
1051 => "001101100",
1052 => "001101101",
1053 => "001101011",
1054 => "001101010",
1055 => "001101001",
1056 => "001101001",
1057 => "001101000",
1058 => "001100111",
1059 => "001101001",
1060 => "001101100",
1061 => "001101001",
1062 => "001101000",
1063 => "001101100",
1064 => "001101011",
1065 => "001101010",
1066 => "001100110",
1067 => "001101000",
1068 => "001100111",
1069 => "001100100",
1070 => "001100110",
1071 => "001100111",
1072 => "001100110",
1073 => "001100101",
1074 => "001100101",
1075 => "001100101",
1076 => "001100110",
1077 => "001100101",
1078 => "001101011",
1079 => "001101100",
1080 => "001101101",
1081 => "001101100",
1082 => "001101101",
1083 => "001101111",
1084 => "001101110",
1085 => "001101111",
1086 => "001101101",
1087 => "001110001",
1088 => "001110000",
1089 => "001110001",
1090 => "001110000",
1091 => "001101011",
1092 => "001101011",
1093 => "001101000",
1094 => "001101010",
1095 => "001101000",
1096 => "001100110",
1097 => "001100110",
1098 => "001100110",
1099 => "001101000",
1100 => "001100101",
1101 => "001101000",
1102 => "001101010",
1103 => "001101000",
1104 => "001101010",
1105 => "001101101",
1106 => "001101111",
1107 => "001101111",
1108 => "001101110",
1109 => "001101010",
1110 => "001101101",
1111 => "001101011",
1112 => "001011100",
1113 => "001010101",
1114 => "001010100",
1115 => "001100001",
1116 => "001101100",
1117 => "001101100",
1118 => "001101010",
1119 => "001101000",
1120 => "001101000",
1121 => "001101100",
1122 => "001101101",
1123 => "001101101",
1124 => "001110000",
1125 => "001110101",
1126 => "001110100",
1127 => "001110101",
1128 => "001110101",
1129 => "001101100",
1130 => "001101011",
1131 => "001101100",
1132 => "001101001",
1133 => "001101011",
1134 => "001101010",
1135 => "001101001",
1136 => "001101111",
1137 => "001101000",
1138 => "001101111",
1139 => "001101011",
1140 => "001101101",
1141 => "001101001",
1142 => "001100111",
1143 => "001101100",
1144 => "001100010",
1145 => "001100010",
1146 => "001100111",
1147 => "001100100",
1148 => "001101000",
1149 => "001100100",
1150 => "001100001",
1151 => "001100110",
1152 => "001100101",
1153 => "001100110",
1154 => "001100101",
1155 => "001011111",
1156 => "001101001",
1157 => "001101001",
1158 => "001101100",
1159 => "001101010",
1160 => "001101110",
1161 => "001101100",
1162 => "001101011",
1163 => "001101001",
1164 => "001101001",
1165 => "001101010",
1166 => "001101100",
1167 => "001100100",
1168 => "001101001",
1169 => "001101100",
1170 => "001101001",
1171 => "001101001",
1172 => "001101011",
1173 => "001101001",
1174 => "001101000",
1175 => "001101001",
1176 => "001100110",
1177 => "001100111",
1178 => "001101010",
1179 => "001101000",
1180 => "001100110",
1181 => "001101010",
1182 => "001100110",
1183 => "001101000",
1184 => "001101001",
1185 => "001101011",
1186 => "001101100",
1187 => "001101100",
1188 => "001101001",
1189 => "001101000",
1190 => "001101001",
1191 => "001101000",
1192 => "001101010",
1193 => "001101001",
1194 => "001100111",
1195 => "001100101",
1196 => "001100011",
1197 => "001100111",
1198 => "001100110",
1199 => "001100100",
1200 => "001100011",
1201 => "001100110",
1202 => "001100101",
1203 => "001100101",
1204 => "001100100",
1205 => "001100011",
1206 => "001100100",
1207 => "001100111",
1208 => "001101000",
1209 => "001100111",
1210 => "001101010",
1211 => "001101101",
1212 => "001101111",
1213 => "001101110",
1214 => "001101000",
1215 => "001101011",
1216 => "001101011",
1217 => "001101101",
1218 => "001101101",
1219 => "001110000",
1220 => "001101110",
1221 => "001101001",
1222 => "001100111",
1223 => "001100111",
1224 => "001101010",
1225 => "001100111",
1226 => "001100111",
1227 => "001100110",
1228 => "001101011",
1229 => "001101010",
1230 => "001101010",
1231 => "001101001",
1232 => "001101100",
1233 => "001101111",
1234 => "001101000",
1235 => "001010011",
1236 => "001100000",
1237 => "001101100",
1238 => "001101011",
1239 => "001100001",
1240 => "001010011",
1241 => "001011000",
1242 => "001011011",
1243 => "001010110",
1244 => "001100010",
1245 => "001100111",
1246 => "001110010",
1247 => "001101110",
1248 => "001110010",
1249 => "001110011",
1250 => "001110101",
1251 => "001101111",
1252 => "001101101",
1253 => "001101001",
1254 => "001110000",
1255 => "001101011",
1256 => "001101001",
1257 => "001101100",
1258 => "001100101",
1259 => "001101110",
1260 => "001101101",
1261 => "001101101",
1262 => "001101011",
1263 => "001101010",
1264 => "001101110",
1265 => "001101101",
1266 => "001101100",
1267 => "001101101",
1268 => "001101010",
1269 => "001101001",
1270 => "001100111",
1271 => "001101000",
1272 => "001100010",
1273 => "001100011",
1274 => "001100110",
1275 => "001100000",
1276 => "001100000",
1277 => "001100010",
1278 => "001100011",
1279 => "001100011",
1280 => "001101000",
1281 => "001100110",
1282 => "001100011",
1283 => "001100100",
1284 => "001101001",
1285 => "001101001",
1286 => "001101011",
1287 => "001101010",
1288 => "001101010",
1289 => "001100100",
1290 => "001100111",
1291 => "001100101",
1292 => "001100110",
1293 => "001101000",
1294 => "001101000",
1295 => "001100111",
1296 => "001101001",
1297 => "001100101",
1298 => "001100111",
1299 => "001100100",
1300 => "001100111",
1301 => "001101000",
1302 => "001100110",
1303 => "001100110",
1304 => "001100111",
1305 => "001100110",
1306 => "001100011",
1307 => "001100101",
1308 => "001100011",
1309 => "001100110",
1310 => "001100110",
1311 => "001100110",
1312 => "001100110",
1313 => "001100101",
1314 => "001100111",
1315 => "001100111",
1316 => "001100100",
1317 => "001100110",
1318 => "001101000",
1319 => "001100111",
1320 => "001101000",
1321 => "001101000",
1322 => "001101001",
1323 => "001101011",
1324 => "001101001",
1325 => "001101010",
1326 => "001101001",
1327 => "001101000",
1328 => "001101010",
1329 => "001101011",
1330 => "001101100",
1331 => "001100101",
1332 => "001100100",
1333 => "001100011",
1334 => "001100100",
1335 => "001100101",
1336 => "001100110",
1337 => "001100111",
1338 => "001101010",
1339 => "001101001",
1340 => "001100110",
1341 => "001101000",
1342 => "001101101",
1343 => "001101110",
1344 => "001101100",
1345 => "001101111",
1346 => "001110000",
1347 => "001110000",
1348 => "001101111",
1349 => "001101011",
1350 => "001101001",
1351 => "001101101",
1352 => "001101010",
1353 => "001101001",
1354 => "001101011",
1355 => "001101001",
1356 => "001100111",
1357 => "001101100",
1358 => "001101100",
1359 => "001101011",
1360 => "001100110",
1361 => "001010100",
1362 => "001010011",
1363 => "001010010",
1364 => "001011101",
1365 => "001101100",
1366 => "001101101",
1367 => "001000100",
1368 => "001000001",
1369 => "001010001",
1370 => "001010000",
1371 => "001110110",
1372 => "001110011",
1373 => "001110111",
1374 => "001111001",
1375 => "001111010",
1376 => "001110011",
1377 => "001101001",
1378 => "001100110",
1379 => "001101111",
1380 => "001101010",
1381 => "001101110",
1382 => "001101100",
1383 => "001101111",
1384 => "001110000",
1385 => "001101111",
1386 => "001100110",
1387 => "001101101",
1388 => "001101101",
1389 => "001110001",
1390 => "001101101",
1391 => "001101011",
1392 => "001101101",
1393 => "001101001",
1394 => "001101111",
1395 => "001101010",
1396 => "001100111",
1397 => "001100011",
1398 => "001100101",
1399 => "001100001",
1400 => "001100110",
1401 => "001100100",
1402 => "001100101",
1403 => "001100100",
1404 => "001100001",
1405 => "001100010",
1406 => "001100100",
1407 => "001011111",
1408 => "001011101",
1409 => "001100100",
1410 => "001100011",
1411 => "001100011",
1412 => "001100111",
1413 => "001100110",
1414 => "001101000",
1415 => "001100111",
1416 => "001101001",
1417 => "001101010",
1418 => "001101000",
1419 => "001101001",
1420 => "001100101",
1421 => "001100110",
1422 => "001101000",
1423 => "001101001",
1424 => "001101101",
1425 => "001101011",
1426 => "001101011",
1427 => "001101011",
1428 => "001101010",
1429 => "001101011",
1430 => "001101010",
1431 => "001100111",
1432 => "001101000",
1433 => "001101000",
1434 => "001100100",
1435 => "001100111",
1436 => "001100101",
1437 => "001011111",
1438 => "001100100",
1439 => "001100110",
1440 => "001101000",
1441 => "001100111",
1442 => "001101010",
1443 => "001101001",
1444 => "001100100",
1445 => "001100111",
1446 => "001100101",
1447 => "001101001",
1448 => "001101000",
1449 => "001101001",
1450 => "001101010",
1451 => "001101001",
1452 => "001101101",
1453 => "001110001",
1454 => "001110011",
1455 => "001110011",
1456 => "001101111",
1457 => "001101101",
1458 => "001101110",
1459 => "001101110",
1460 => "001101101",
1461 => "001101111",
1462 => "001101001",
1463 => "001101101",
1464 => "001101110",
1465 => "001101111",
1466 => "001101100",
1467 => "001101111",
1468 => "001101110",
1469 => "001110010",
1470 => "001110010",
1471 => "001110001",
1472 => "001110001",
1473 => "001101111",
1474 => "001101110",
1475 => "001101111",
1476 => "001101111",
1477 => "001101110",
1478 => "001101001",
1479 => "001101001",
1480 => "001101100",
1481 => "001101110",
1482 => "001101111",
1483 => "001101111",
1484 => "001110000",
1485 => "001101111",
1486 => "001110000",
1487 => "001011110",
1488 => "001010110",
1489 => "001010101",
1490 => "001011001",
1491 => "001010111",
1492 => "001011010",
1493 => "001101100",
1494 => "001101101",
1495 => "001011011",
1496 => "001010111",
1497 => "001101001",
1498 => "001101001",
1499 => "001110000",
1500 => "001101011",
1501 => "001101000",
1502 => "001100111",
1503 => "001110001",
1504 => "001101111",
1505 => "001101110",
1506 => "001101101",
1507 => "001101010",
1508 => "001110000",
1509 => "001110011",
1510 => "001110100",
1511 => "001110011",
1512 => "001110010",
1513 => "001110011",
1514 => "001101100",
1515 => "001101110",
1516 => "001101110",
1517 => "001110000",
1518 => "001101011",
1519 => "001110000",
1520 => "001110000",
1521 => "001101111",
1522 => "001101111",
1523 => "001101001",
1524 => "001101011",
1525 => "001100101",
1526 => "001100111",
1527 => "001100110",
1528 => "001100110",
1529 => "001100100",
1530 => "001100100",
1531 => "001100100",
1532 => "001100011",
1533 => "001100001",
1534 => "001100010",
1535 => "001100010",
1536 => "001101000",
1537 => "001100111",
1538 => "001100101",
1539 => "001100011",
1540 => "001100011",
1541 => "001100101",
1542 => "001101000",
1543 => "001101010",
1544 => "001101010",
1545 => "001101011",
1546 => "001101000",
1547 => "001100011",
1548 => "001100111",
1549 => "001100100",
1550 => "001100100",
1551 => "001101000",
1552 => "001101001",
1553 => "001101010",
1554 => "001101010",
1555 => "001100100",
1556 => "001101011",
1557 => "001101010",
1558 => "001101001",
1559 => "001101001",
1560 => "001101000",
1561 => "001100101",
1562 => "001100011",
1563 => "001100101",
1564 => "001100011",
1565 => "001100101",
1566 => "001100010",
1567 => "001100101",
1568 => "001100101",
1569 => "001100111",
1570 => "001101000",
1571 => "001101011",
1572 => "001101001",
1573 => "001101111",
1574 => "001101101",
1575 => "001101101",
1576 => "001101101",
1577 => "001101101",
1578 => "001101101",
1579 => "001101101",
1580 => "001110000",
1581 => "001111001",
1582 => "001110101",
1583 => "001100101",
1584 => "001101011",
1585 => "001101011",
1586 => "001101100",
1587 => "001101100",
1588 => "001101100",
1589 => "001101100",
1590 => "001101110",
1591 => "001101101",
1592 => "001101011",
1593 => "001101010",
1594 => "001101010",
1595 => "001101011",
1596 => "001110000",
1597 => "001101101",
1598 => "001101100",
1599 => "001101100",
1600 => "001110000",
1601 => "001110000",
1602 => "001101110",
1603 => "001101111",
1604 => "001110000",
1605 => "001110001",
1606 => "001110000",
1607 => "001110000",
1608 => "001101111",
1609 => "001110011",
1610 => "001111010",
1611 => "001110101",
1612 => "001111001",
1613 => "001110111",
1614 => "001110100",
1615 => "001110100",
1616 => "001110110",
1617 => "001101100",
1618 => "001101100",
1619 => "001110010",
1620 => "001110010",
1621 => "001110000",
1622 => "001110001",
1623 => "001110001",
1624 => "001110000",
1625 => "001110001",
1626 => "001101111",
1627 => "001101110",
1628 => "001110011",
1629 => "001110111",
1630 => "001110101",
1631 => "001110011",
1632 => "001110011",
1633 => "001110000",
1634 => "001110100",
1635 => "001110011",
1636 => "001110011",
1637 => "001101100",
1638 => "001110000",
1639 => "001110001",
1640 => "001101111",
1641 => "001101101",
1642 => "001101101",
1643 => "001101111",
1644 => "001101101",
1645 => "001101110",
1646 => "001101001",
1647 => "001101000",
1648 => "001101010",
1649 => "001101010",
1650 => "001100010",
1651 => "001100001",
1652 => "001100010",
1653 => "001011101",
1654 => "001100011",
1655 => "001100011",
1656 => "001100111",
1657 => "001101001",
1658 => "001100111",
1659 => "001100100",
1660 => "001100011",
1661 => "001011110",
1662 => "001011100",
1663 => "001100000",
1664 => "001100100",
1665 => "001100111",
1666 => "001101001",
1667 => "001101000",
1668 => "001100111",
1669 => "001101010",
1670 => "001100111",
1671 => "001101000",
1672 => "001100010",
1673 => "001100100",
1674 => "001100100",
1675 => "001100101",
1676 => "001100010",
1677 => "001100111",
1678 => "001100111",
1679 => "001100110",
1680 => "001100110",
1681 => "001100101",
1682 => "001101001",
1683 => "001100101",
1684 => "001100101",
1685 => "001101000",
1686 => "001101001",
1687 => "001101001",
1688 => "001100100",
1689 => "001100111",
1690 => "001101001",
1691 => "001100111",
1692 => "001100011",
1693 => "001101000",
1694 => "001101000",
1695 => "001101001",
1696 => "001101010",
1697 => "001100011",
1698 => "001100111",
1699 => "001101000",
1700 => "001101100",
1701 => "001101010",
1702 => "001101100",
1703 => "001101010",
1704 => "001101000",
1705 => "001101011",
1706 => "001101011",
1707 => "001110001",
1708 => "001101100",
1709 => "001100110",
1710 => "001100100",
1711 => "001100001",
1712 => "001101100",
1713 => "001101110",
1714 => "001101011",
1715 => "001101010",
1716 => "001101010",
1717 => "001101100",
1718 => "001101001",
1719 => "001101000",
1720 => "001101011",
1721 => "001100111",
1722 => "001101001",
1723 => "001100101",
1724 => "001101011",
1725 => "001100100",
1726 => "001101001",
1727 => "001101010",
1728 => "001101110",
1729 => "001110101",
1730 => "001110100",
1731 => "001110110",
1732 => "001111000",
1733 => "001110101",
1734 => "001110011",
1735 => "001110011",
1736 => "001101110",
1737 => "001110010",
1738 => "001110111",
1739 => "001110011",
1740 => "001101001",
1741 => "001101010",
1742 => "001101011",
1743 => "001101110",
1744 => "001101111",
1745 => "001110001",
1746 => "001101101",
1747 => "001101010",
1748 => "001101011",
1749 => "001101001",
1750 => "001101000",
1751 => "001101101",
1752 => "001101011",
1753 => "001110000",
1754 => "001101100",
1755 => "001101000",
1756 => "001100111",
1757 => "001101010",
1758 => "001110010",
1759 => "001101111",
1760 => "001101101",
1761 => "001101100",
1762 => "001101101",
1763 => "001101101",
1764 => "001101010",
1765 => "001101011",
1766 => "001101001",
1767 => "001101001",
1768 => "001101011",
1769 => "001100111",
1770 => "001101001",
1771 => "001100101",
1772 => "001100101",
1773 => "001100101",
1774 => "001100011",
1775 => "001100101",
1776 => "001101000",
1777 => "001100100",
1778 => "001100111",
1779 => "001101010",
1780 => "001101011",
1781 => "001101001",
1782 => "001101011",
1783 => "001101010",
1784 => "001100110",
1785 => "001100110",
1786 => "001100111",
1787 => "001100110",
1788 => "001100111",
1789 => "001100111",
1790 => "001011111",
1791 => "001100010",
1792 => "001100100",
1793 => "001100011",
1794 => "001100011",
1795 => "001100000",
1796 => "001100010",
1797 => "001100000",
1798 => "001011110",
1799 => "001100000",
1800 => "001100010",
1801 => "001100100",
1802 => "001011010",
1803 => "001100001",
1804 => "001011111",
1805 => "001100101",
1806 => "001100000",
1807 => "001100100",
1808 => "001100001",
1809 => "001100101",
1810 => "001011111",
1811 => "001100110",
1812 => "001100011",
1813 => "001100110",
1814 => "001100010",
1815 => "001100011",
1816 => "001100110",
1817 => "001100011",
1818 => "001100011",
1819 => "001100100",
1820 => "001100011",
1821 => "001100101",
1822 => "001101001",
1823 => "001100101",
1824 => "001100100",
1825 => "001100100",
1826 => "001101000",
1827 => "001100101",
1828 => "001100101",
1829 => "001101000",
1830 => "001100101",
1831 => "001101001",
1832 => "001101011",
1833 => "001101010",
1834 => "001101100",
1835 => "001101000",
1836 => "001101001",
1837 => "001101100",
1838 => "001100110",
1839 => "001101110",
1840 => "001110011",
1841 => "001101111",
1842 => "001101111",
1843 => "001101110",
1844 => "001101100",
1845 => "001101001",
1846 => "001101110",
1847 => "001101100",
1848 => "001101001",
1849 => "001101001",
1850 => "001100110",
1851 => "001100111",
1852 => "001101011",
1853 => "001101110",
1854 => "001110011",
1855 => "001101111",
1856 => "001101110",
1857 => "001110010",
1858 => "001110001",
1859 => "001101100",
1860 => "001101100",
1861 => "001101101",
1862 => "001101111",
1863 => "001110010",
1864 => "001101101",
1865 => "001101010",
1866 => "001101010",
1867 => "001101110",
1868 => "001101100",
1869 => "001101010",
1870 => "001110000",
1871 => "001101110",
1872 => "001101011",
1873 => "001101111",
1874 => "001110000",
1875 => "001101001",
1876 => "001101110",
1877 => "001101011",
1878 => "001101101",
1879 => "001101110",
1880 => "001101100",
1881 => "001110000",
1882 => "001101101",
1883 => "001101111",
1884 => "001101110",
1885 => "001101100",
1886 => "001101111",
1887 => "001101110",
1888 => "001101111",
1889 => "001101100",
1890 => "001101100",
1891 => "001101011",
1892 => "001101100",
1893 => "001101111",
1894 => "001101010",
1895 => "001101000",
1896 => "001101101",
1897 => "001101011",
1898 => "001101011",
1899 => "001101110",
1900 => "001101000",
1901 => "001100100",
1902 => "001101011",
1903 => "001101001",
1904 => "001101100",
1905 => "001101101",
1906 => "001101101",
1907 => "001101010",
1908 => "001101101",
1909 => "001100111",
1910 => "001100101",
1911 => "001100100",
1912 => "001100000",
1913 => "001100001",
1914 => "001100011",
1915 => "001100100",
1916 => "001100001",
1917 => "001100111",
1918 => "001100000",
1919 => "001011100",
1920 => "001100101",
1921 => "001100100",
1922 => "001100110",
1923 => "001100101",
1924 => "001100001",
1925 => "001100100",
1926 => "001011100",
1927 => "001100110",
1928 => "001100010",
1929 => "001011001",
1930 => "001011101",
1931 => "001011111",
1932 => "001100010",
1933 => "001100000",
1934 => "001100001",
1935 => "001100010",
1936 => "001100010",
1937 => "001100010",
1938 => "001100001",
1939 => "001100100",
1940 => "001100100",
1941 => "001100010",
1942 => "001100011",
1943 => "001100011",
1944 => "001100001",
1945 => "001100110",
1946 => "001100011",
1947 => "001100000",
1948 => "001100001",
1949 => "001011110",
1950 => "001100010",
1951 => "001100100",
1952 => "001100001",
1953 => "001100010",
1954 => "001100010",
1955 => "001011111",
1956 => "001100010",
1957 => "001100001",
1958 => "001100011",
1959 => "001100101",
1960 => "001100011",
1961 => "001100011",
1962 => "001100011",
1963 => "001011110",
1964 => "001100100",
1965 => "001101000",
1966 => "001011100",
1967 => "001010100",
1968 => "001100000",
1969 => "001100011",
1970 => "001101011",
1971 => "001101001",
1972 => "001100010",
1973 => "001101100",
1974 => "001101011",
1975 => "001101100",
1976 => "001101001",
1977 => "001110000",
1978 => "001110010",
1979 => "001110111",
1980 => "001101110",
1981 => "001101110",
1982 => "001101111",
1983 => "001101100",
1984 => "001101111",
1985 => "001101001",
1986 => "001101011",
1987 => "001101010",
1988 => "001110001",
1989 => "001101111",
1990 => "001101100",
1991 => "001101100",
1992 => "001101100",
1993 => "001110011",
1994 => "001101100",
1995 => "001101010",
1996 => "001101101",
1997 => "001101100",
1998 => "001101110",
1999 => "001100110",
2000 => "001101011",
2001 => "001101010",
2002 => "001101010",
2003 => "001101100",
2004 => "001101011",
2005 => "001101100",
2006 => "001101100",
2007 => "001101001",
2008 => "001101010",
2009 => "001101010",
2010 => "001101011",
2011 => "001101010",
2012 => "001101100",
2013 => "001101000",
2014 => "001101101",
2015 => "001101001",
2016 => "001101010",
2017 => "001101100",
2018 => "001101010",
2019 => "001101010",
2020 => "001101011",
2021 => "001101100",
2022 => "001110000",
2023 => "001110000",
2024 => "001101101",
2025 => "001101101",
2026 => "001101101",
2027 => "001101110",
2028 => "001101011",
2029 => "001101000",
2030 => "001101100",
2031 => "001100111",
2032 => "001100001",
2033 => "001100101",
2034 => "001100111",
2035 => "001100000",
2036 => "001100101",
2037 => "001100011",
2038 => "001100111",
2039 => "001100001",
2040 => "001100000",
2041 => "001011100",
2042 => "001011111",
2043 => "001011111",
2044 => "001011101",
2045 => "001011101",
2046 => "001011110",
2047 => "001011101",
2048 => "001100001",
2049 => "001100111",
2050 => "001100011",
2051 => "001100010",
2052 => "001100001",
2053 => "001100011",
2054 => "001011101",
2055 => "001100001",
2056 => "001010100",
2057 => "001011100",
2058 => "001100001",
2059 => "001011111",
2060 => "001011101",
2061 => "001100101",
2062 => "001100011",
2063 => "001100001",
2064 => "001100010",
2065 => "001100001",
2066 => "001100101",
2067 => "001100101",
2068 => "001100010",
2069 => "001100010",
2070 => "001100000",
2071 => "001100000",
2072 => "001100100",
2073 => "001100000",
2074 => "001100010",
2075 => "001100011",
2076 => "001100110",
2077 => "001011111",
2078 => "001100001",
2079 => "001100001",
2080 => "001100010",
2081 => "001011111",
2082 => "001100010",
2083 => "001100101",
2084 => "001100011",
2085 => "001101010",
2086 => "001101101",
2087 => "001101100",
2088 => "001100101",
2089 => "001100110",
2090 => "001101000",
2091 => "001100001",
2092 => "001101100",
2093 => "001101111",
2094 => "001100111",
2095 => "001101100",
2096 => "001101011",
2097 => "001100111",
2098 => "001101001",
2099 => "001101111",
2100 => "001100111",
2101 => "001101001",
2102 => "001101101",
2103 => "001110010",
2104 => "001110011",
2105 => "001110001",
2106 => "001110101",
2107 => "001101111",
2108 => "001110011",
2109 => "001110000",
2110 => "001110011",
2111 => "001101111",
2112 => "001110001",
2113 => "001101111",
2114 => "001110001",
2115 => "001101101",
2116 => "001101110",
2117 => "001101111",
2118 => "001110001",
2119 => "001101111",
2120 => "001110001",
2121 => "001101101",
2122 => "001101110",
2123 => "001101110",
2124 => "001101101",
2125 => "001101110",
2126 => "001101100",
2127 => "001101101",
2128 => "001101111",
2129 => "001101110",
2130 => "001101011",
2131 => "001101010",
2132 => "001101011",
2133 => "001101000",
2134 => "001101000",
2135 => "001101000",
2136 => "001101011",
2137 => "001101100",
2138 => "001101010",
2139 => "001101000",
2140 => "001101111",
2141 => "001101010",
2142 => "001101010",
2143 => "001101000",
2144 => "001101011",
2145 => "001101110",
2146 => "001101110",
2147 => "001101001",
2148 => "001101111",
2149 => "001101101",
2150 => "001101100",
2151 => "001101011",
2152 => "001100101",
2153 => "001100111",
2154 => "001101100",
2155 => "001101110",
2156 => "001101010",
2157 => "001101010",
2158 => "001101100",
2159 => "001100111",
2160 => "001101000",
2161 => "001100111",
2162 => "001100111",
2163 => "001101001",
2164 => "001100110",
2165 => "001100110",
2166 => "001100100",
2167 => "001100111",
2168 => "001101000",
2169 => "001101000",
2170 => "001100011",
2171 => "001100001",
2172 => "001100001",
2173 => "001100001",
2174 => "001100000",
2175 => "001100001",
2176 => "001100001",
2177 => "001100001",
2178 => "001100000",
2179 => "001100011",
2180 => "001100101",
2181 => "001100100",
2182 => "001100010",
2183 => "001100001",
2184 => "001100011",
2185 => "001100011",
2186 => "001011111",
2187 => "001100101",
2188 => "001100010",
2189 => "001100010",
2190 => "001100001",
2191 => "001011100",
2192 => "001011111",
2193 => "001100011",
2194 => "001100100",
2195 => "001100101",
2196 => "001100110",
2197 => "001100010",
2198 => "001011111",
2199 => "001101010",
2200 => "001101000",
2201 => "001101001",
2202 => "001101010",
2203 => "001101001",
2204 => "001101010",
2205 => "001101110",
2206 => "001101010",
2207 => "001101001",
2208 => "001101001",
2209 => "001101101",
2210 => "001011110",
2211 => "001100000",
2212 => "001100011",
2213 => "001011010",
2214 => "001100110",
2215 => "001100100",
2216 => "001011001",
2217 => "001100101",
2218 => "001011101",
2219 => "001101000",
2220 => "001101100",
2221 => "001101111",
2222 => "001101100",
2223 => "001101101",
2224 => "001101100",
2225 => "001101111",
2226 => "001101110",
2227 => "001101110",
2228 => "001110011",
2229 => "001111010",
2230 => "001110101",
2231 => "001111001",
2232 => "001110010",
2233 => "001110011",
2234 => "001110100",
2235 => "001101111",
2236 => "001110001",
2237 => "001110000",
2238 => "001101110",
2239 => "001110000",
2240 => "001101100",
2241 => "001101111",
2242 => "001101111",
2243 => "001101111",
2244 => "001101111",
2245 => "001101101",
2246 => "001101111",
2247 => "001110000",
2248 => "001110011",
2249 => "001110011",
2250 => "001110100",
2251 => "001110000",
2252 => "001110000",
2253 => "001110010",
2254 => "001110010",
2255 => "001110010",
2256 => "001110000",
2257 => "001101100",
2258 => "001101100",
2259 => "001101110",
2260 => "001101111",
2261 => "001101100",
2262 => "001101011",
2263 => "001100101",
2264 => "001101010",
2265 => "001101001",
2266 => "001101010",
2267 => "001101011",
2268 => "001101001",
2269 => "001101100",
2270 => "001101000",
2271 => "001101011",
2272 => "001100101",
2273 => "001101010",
2274 => "001101010",
2275 => "001101000",
2276 => "001100110",
2277 => "001100101",
2278 => "001100111",
2279 => "001110001",
2280 => "001101110",
2281 => "001101001",
2282 => "001101000",
2283 => "001101001",
2284 => "001101010",
2285 => "001101011",
2286 => "001101110",
2287 => "001101001",
2288 => "001101010",
2289 => "001101010",
2290 => "001100111",
2291 => "001101001",
2292 => "001101011",
2293 => "001100111",
2294 => "001100111",
2295 => "001100101",
2296 => "001100010",
2297 => "001100100",
2298 => "001100111",
2299 => "001101000",
2300 => "001100101",
2301 => "001100100",
2302 => "001011111",
2303 => "001011100",
2304 => "001100001",
2305 => "001100110",
2306 => "001011111",
2307 => "001100101",
2308 => "001100111",
2309 => "001101001",
2310 => "001100110",
2311 => "001101000",
2312 => "001100111",
2313 => "001101010",
2314 => "001100101",
2315 => "001100110",
2316 => "001100111",
2317 => "001101010",
2318 => "001101010",
2319 => "001101000",
2320 => "001101110",
2321 => "001101000",
2322 => "001101101",
2323 => "001101100",
2324 => "001101000",
2325 => "001110000",
2326 => "001101001",
2327 => "001101001",
2328 => "001100101",
2329 => "001100011",
2330 => "001100100",
2331 => "001100111",
2332 => "001101011",
2333 => "001101001",
2334 => "001101010",
2335 => "001100011",
2336 => "001011100",
2337 => "001011111",
2338 => "001100100",
2339 => "001011111",
2340 => "001100001",
2341 => "001101111",
2342 => "001101000",
2343 => "001110000",
2344 => "001101111",
2345 => "001101100",
2346 => "001110011",
2347 => "001101111",
2348 => "001110101",
2349 => "001110000",
2350 => "001110011",
2351 => "001110010",
2352 => "001110101",
2353 => "001110100",
2354 => "001110001",
2355 => "001110000",
2356 => "001101111",
2357 => "001101111",
2358 => "001101110",
2359 => "001101101",
2360 => "001110001",
2361 => "001101110",
2362 => "001101111",
2363 => "001101011",
2364 => "001101100",
2365 => "001101100",
2366 => "001101110",
2367 => "001101100",
2368 => "001101101",
2369 => "001101100",
2370 => "001110010",
2371 => "001110001",
2372 => "001101111",
2373 => "001110010",
2374 => "001110010",
2375 => "001101111",
2376 => "001101101",
2377 => "001101111",
2378 => "001101110",
2379 => "001101111",
2380 => "001101101",
2381 => "001110000",
2382 => "001110000",
2383 => "001110011",
2384 => "001110101",
2385 => "001110110",
2386 => "001110011",
2387 => "001110001",
2388 => "001101110",
2389 => "001101111",
2390 => "001101101",
2391 => "001101101",
2392 => "001101011",
2393 => "001100101",
2394 => "001100111",
2395 => "001100010",
2396 => "001100001",
2397 => "001100101",
2398 => "001100111",
2399 => "001101001",
2400 => "001101010",
2401 => "001101101",
2402 => "001101000",
2403 => "001100111",
2404 => "001101001",
2405 => "001100001",
2406 => "001100100",
2407 => "001100101",
2408 => "001100110",
2409 => "001100100",
2410 => "001101000",
2411 => "001101010",
2412 => "001101010",
2413 => "001100111",
2414 => "001100111",
2415 => "001100010",
2416 => "001100101",
2417 => "001100011",
2418 => "001100000",
2419 => "001100001",
2420 => "001100100",
2421 => "001100110",
2422 => "001100100",
2423 => "001100100",
2424 => "001100100",
2425 => "001100010",
2426 => "001011111",
2427 => "001100000",
2428 => "001011000",
2429 => "001011100",
2430 => "001100001",
2431 => "001011101",
2432 => "001110001",
2433 => "001110110",
2434 => "001111010",
2435 => "001110100",
2436 => "001111000",
2437 => "001111011",
2438 => "001110011",
2439 => "001110110",
2440 => "001101111",
2441 => "001100101",
2442 => "001101100",
2443 => "001101000",
2444 => "001100110",
2445 => "001100110",
2446 => "001100001",
2447 => "001100101",
2448 => "001011010",
2449 => "001100000",
2450 => "001100101",
2451 => "001100110",
2452 => "001011111",
2453 => "001101001",
2454 => "001100111",
2455 => "001101000",
2456 => "001011111",
2457 => "001100111",
2458 => "001101000",
2459 => "001100110",
2460 => "001100110",
2461 => "001100111",
2462 => "001011101",
2463 => "001100011",
2464 => "001100100",
2465 => "001101001",
2466 => "001100100",
2467 => "001101011",
2468 => "001101010",
2469 => "001110001",
2470 => "001110000",
2471 => "001101101",
2472 => "001101101",
2473 => "001101110",
2474 => "001101010",
2475 => "001101101",
2476 => "001101100",
2477 => "001110000",
2478 => "001101111",
2479 => "001110001",
2480 => "001101111",
2481 => "001110001",
2482 => "001110000",
2483 => "001110000",
2484 => "001101110",
2485 => "001101011",
2486 => "001101000",
2487 => "001101010",
2488 => "001101001",
2489 => "001101100",
2490 => "001101001",
2491 => "001101011",
2492 => "001101101",
2493 => "001101010",
2494 => "001101010",
2495 => "001101011",
2496 => "001101001",
2497 => "001101110",
2498 => "001101101",
2499 => "001101111",
2500 => "001101011",
2501 => "001110001",
2502 => "001101011",
2503 => "001101100",
2504 => "001101001",
2505 => "001101010",
2506 => "001101011",
2507 => "001101100",
2508 => "001101101",
2509 => "001110001",
2510 => "001101101",
2511 => "001101111",
2512 => "001101101",
2513 => "001101101",
2514 => "001110001",
2515 => "001101010",
2516 => "001101000",
2517 => "001101000",
2518 => "001101011",
2519 => "001101011",
2520 => "001101010",
2521 => "001100101",
2522 => "001101001",
2523 => "001101011",
2524 => "001100111",
2525 => "001100110",
2526 => "001101010",
2527 => "001100110",
2528 => "001101001",
2529 => "001101001",
2530 => "001100111",
2531 => "001100110",
2532 => "001100111",
2533 => "001101010",
2534 => "001101010",
2535 => "001100100",
2536 => "001101010",
2537 => "001101001",
2538 => "001100011",
2539 => "001100100",
2540 => "001100011",
2541 => "001100100",
2542 => "001100110",
2543 => "001100011",
2544 => "001100100",
2545 => "001100110",
2546 => "001100000",
2547 => "001100010",
2548 => "001100001",
2549 => "001011101",
2550 => "001011001",
2551 => "001011110",
2552 => "001100000",
2553 => "001100011",
2554 => "001011011",
2555 => "001100010",
2556 => "001100010",
2557 => "001100011",
2558 => "001100000",
2559 => "001100000",
2560 => "001101100",
2561 => "001101010",
2562 => "001100100",
2563 => "001100110",
2564 => "001101011",
2565 => "001101010",
2566 => "001100111",
2567 => "001101000",
2568 => "001100011",
2569 => "001011100",
2570 => "001011111",
2571 => "001011011",
2572 => "001100010",
2573 => "001011110",
2574 => "001011110",
2575 => "001011100",
2576 => "001011111",
2577 => "001100000",
2578 => "001011100",
2579 => "001100001",
2580 => "001100010",
2581 => "001100010",
2582 => "001100000",
2583 => "001100011",
2584 => "001011001",
2585 => "001011101",
2586 => "001011101",
2587 => "001100001",
2588 => "001011100",
2589 => "001100010",
2590 => "001101010",
2591 => "001110000",
2592 => "001101100",
2593 => "001101101",
2594 => "001100100",
2595 => "001101000",
2596 => "001101110",
2597 => "001101100",
2598 => "001101100",
2599 => "001101011",
2600 => "001101000",
2601 => "001101111",
2602 => "001101111",
2603 => "001101111",
2604 => "001101111",
2605 => "001110001",
2606 => "001101010",
2607 => "001101101",
2608 => "001101101",
2609 => "001101101",
2610 => "001101101",
2611 => "001100111",
2612 => "001101010",
2613 => "001101000",
2614 => "001100111",
2615 => "001101011",
2616 => "001100110",
2617 => "001101100",
2618 => "001101001",
2619 => "001100101",
2620 => "001101100",
2621 => "001100111",
2622 => "001101100",
2623 => "001101000",
2624 => "001101000",
2625 => "001101001",
2626 => "001101111",
2627 => "001101011",
2628 => "001101000",
2629 => "001101101",
2630 => "001101101",
2631 => "001101011",
2632 => "001101010",
2633 => "001101001",
2634 => "001101010",
2635 => "001101100",
2636 => "001101101",
2637 => "001100110",
2638 => "001101011",
2639 => "001101000",
2640 => "001100111",
2641 => "001100101",
2642 => "001100111",
2643 => "001100101",
2644 => "001100100",
2645 => "001100111",
2646 => "001101010",
2647 => "001100111",
2648 => "001101010",
2649 => "001101010",
2650 => "001101011",
2651 => "001101100",
2652 => "001101110",
2653 => "001101110",
2654 => "001101010",
2655 => "001101000",
2656 => "001101000",
2657 => "001101011",
2658 => "001101000",
2659 => "001101001",
2660 => "001101101",
2661 => "001101010",
2662 => "001101011",
2663 => "001100101",
2664 => "001100110",
2665 => "001100101",
2666 => "001100011",
2667 => "001100111",
2668 => "001100111",
2669 => "001100100",
2670 => "001101010",
2671 => "001100100",
2672 => "001100000",
2673 => "001100110",
2674 => "001100010",
2675 => "001100101",
2676 => "001100110",
2677 => "001100010",
2678 => "001100000",
2679 => "001011101",
2680 => "001100010",
2681 => "001010011",
2682 => "001100000",
2683 => "001010110",
2684 => "001011011",
2685 => "001011101",
2686 => "001100000",
2687 => "001011011",
2688 => "001101000",
2689 => "001101001",
2690 => "001101001",
2691 => "001101100",
2692 => "001101011",
2693 => "001101100",
2694 => "001110001",
2695 => "001101000",
2696 => "001011110",
2697 => "001011110",
2698 => "001010111",
2699 => "001011111",
2700 => "001100010",
2701 => "001011111",
2702 => "001100001",
2703 => "001100101",
2704 => "001100100",
2705 => "001101011",
2706 => "001100100",
2707 => "001101000",
2708 => "001100111",
2709 => "001100011",
2710 => "001101110",
2711 => "001101010",
2712 => "001101010",
2713 => "001111000",
2714 => "001110111",
2715 => "001110011",
2716 => "001111101",
2717 => "001111001",
2718 => "001110101",
2719 => "001110001",
2720 => "001110100",
2721 => "001110001",
2722 => "001101101",
2723 => "001101010",
2724 => "001101000",
2725 => "001101111",
2726 => "001101100",
2727 => "001110001",
2728 => "001101100",
2729 => "001110001",
2730 => "001110001",
2731 => "001110001",
2732 => "001101001",
2733 => "001110001",
2734 => "001110001",
2735 => "001101100",
2736 => "001110011",
2737 => "001101000",
2738 => "001101101",
2739 => "001101011",
2740 => "001110010",
2741 => "001100111",
2742 => "001100010",
2743 => "001101001",
2744 => "001101001",
2745 => "001101001",
2746 => "001101010",
2747 => "001101101",
2748 => "001100111",
2749 => "001101001",
2750 => "001101010",
2751 => "001100111",
2752 => "001100111",
2753 => "001100100",
2754 => "001100100",
2755 => "001101001",
2756 => "001101000",
2757 => "001100111",
2758 => "001101011",
2759 => "001101010",
2760 => "001101100",
2761 => "001100101",
2762 => "001100000",
2763 => "001100110",
2764 => "001100101",
2765 => "001100111",
2766 => "001011110",
2767 => "001100011",
2768 => "001100011",
2769 => "001101000",
2770 => "001100000",
2771 => "001101000",
2772 => "001101000",
2773 => "001101000",
2774 => "001100111",
2775 => "001101110",
2776 => "001101000",
2777 => "001100111",
2778 => "001100110",
2779 => "001100111",
2780 => "001100100",
2781 => "001100101",
2782 => "001100010",
2783 => "001100110",
2784 => "001100100",
2785 => "001100011",
2786 => "001100111",
2787 => "001100111",
2788 => "001101000",
2789 => "001100111",
2790 => "001101011",
2791 => "001100111",
2792 => "001100110",
2793 => "001100111",
2794 => "001100010",
2795 => "001100110",
2796 => "001100100",
2797 => "001101000",
2798 => "001101011",
2799 => "001100011",
2800 => "001100011",
2801 => "001110011",
2802 => "001101111",
2803 => "001100110",
2804 => "001100001",
2805 => "001100011",
2806 => "001100011",
2807 => "001100000",
2808 => "001011111",
2809 => "001011111",
2810 => "001011111",
2811 => "001011110",
2812 => "001010100",
2813 => "001011100",
2814 => "001011110",
2815 => "001011000",
2816 => "001011001",
2817 => "001100001",
2818 => "001101000",
2819 => "001101110",
2820 => "001100000",
2821 => "001100000",
2822 => "001100001",
2823 => "001100011",
2824 => "001100000",
2825 => "001011011",
2826 => "001100111",
2827 => "001100010",
2828 => "001011110",
2829 => "001101110",
2830 => "001110011",
2831 => "001101100",
2832 => "001101100",
2833 => "001100000",
2834 => "001100110",
2835 => "001110111",
2836 => "001101110",
2837 => "001110011",
2838 => "001110001",
2839 => "001101011",
2840 => "001101001",
2841 => "001101000",
2842 => "001101100",
2843 => "001101011",
2844 => "001101100",
2845 => "001101100",
2846 => "001101001",
2847 => "001101111",
2848 => "001101000",
2849 => "001101001",
2850 => "001101110",
2851 => "001110010",
2852 => "001101110",
2853 => "001110100",
2854 => "001110001",
2855 => "001110001",
2856 => "001110010",
2857 => "001101110",
2858 => "001101111",
2859 => "001110010",
2860 => "001110011",
2861 => "001110100",
2862 => "001101001",
2863 => "001101100",
2864 => "001110010",
2865 => "001101010",
2866 => "001101101",
2867 => "001101111",
2868 => "001101000",
2869 => "001101000",
2870 => "001110000",
2871 => "001110000",
2872 => "001101001",
2873 => "001100001",
2874 => "001100101",
2875 => "001100110",
2876 => "001101001",
2877 => "001100011",
2878 => "001101000",
2879 => "001100111",
2880 => "001100101",
2881 => "001101001",
2882 => "001100111",
2883 => "001101000",
2884 => "001101000",
2885 => "001100110",
2886 => "001100010",
2887 => "001101101",
2888 => "001100100",
2889 => "001100101",
2890 => "001100001",
2891 => "001111010",
2892 => "001100110",
2893 => "001100000",
2894 => "001100001",
2895 => "001100010",
2896 => "001100100",
2897 => "001101000",
2898 => "001100000",
2899 => "001100011",
2900 => "001101000",
2901 => "001100001",
2902 => "001101100",
2903 => "001101111",
2904 => "001100110",
2905 => "001100100",
2906 => "001101001",
2907 => "001100101",
2908 => "001100000",
2909 => "001100011",
2910 => "001100101",
2911 => "001100111",
2912 => "001100101",
2913 => "001101010",
2914 => "001100110",
2915 => "001101000",
2916 => "001100111",
2917 => "001101010",
2918 => "001110000",
2919 => "001101000",
2920 => "001100100",
2921 => "001101000",
2922 => "001100111",
2923 => "001011101",
2924 => "001011100",
2925 => "001011001",
2926 => "001100001",
2927 => "001100001",
2928 => "001001101",
2929 => "001001011",
2930 => "001011011",
2931 => "001011101",
2932 => "001100111",
2933 => "001100100",
2934 => "001100000",
2935 => "001100100",
2936 => "001100111",
2937 => "001100001",
2938 => "001011011",
2939 => "001100000",
2940 => "001100011",
2941 => "001011100",
2942 => "001100010",
2943 => "001100100",
2944 => "001011001",
2945 => "001010100",
2946 => "001011011",
2947 => "001011110",
2948 => "001101001",
2949 => "001100010",
2950 => "001011111",
2951 => "001100110",
2952 => "001101000",
2953 => "001100110",
2954 => "001101111",
2955 => "001110011",
2956 => "001110000",
2957 => "001110000",
2958 => "001110011",
2959 => "001110000",
2960 => "001110001",
2961 => "001110000",
2962 => "001101111",
2963 => "001110000",
2964 => "001110000",
2965 => "001110000",
2966 => "001110001",
2967 => "001101111",
2968 => "001101111",
2969 => "001101100",
2970 => "001101101",
2971 => "001110101",
2972 => "001101111",
2973 => "001110000",
2974 => "001110000",
2975 => "001110101",
2976 => "001110101",
2977 => "001110011",
2978 => "001110000",
2979 => "001101100",
2980 => "001110010",
2981 => "001101110",
2982 => "001111000",
2983 => "001110001",
2984 => "001101010",
2985 => "001110011",
2986 => "001101101",
2987 => "001100111",
2988 => "001110010",
2989 => "001110000",
2990 => "001110001",
2991 => "001110001",
2992 => "001101110",
2993 => "001101111",
2994 => "001101100",
2995 => "001101111",
2996 => "001101111",
2997 => "001110000",
2998 => "001101010",
2999 => "001101011",
3000 => "001101110",
3001 => "001101111",
3002 => "001101100",
3003 => "001101101",
3004 => "001101011",
3005 => "001101010",
3006 => "001110001",
3007 => "001101010",
3008 => "001101111",
3009 => "001101011",
3010 => "001101001",
3011 => "001101101",
3012 => "001101111",
3013 => "001110011",
3014 => "001101010",
3015 => "001101001",
3016 => "001110011",
3017 => "001101110",
3018 => "001110011",
3019 => "001110000",
3020 => "001101010",
3021 => "001101000",
3022 => "001100011",
3023 => "001110001",
3024 => "001100101",
3025 => "001100110",
3026 => "001011100",
3027 => "001100110",
3028 => "001101100",
3029 => "001100110",
3030 => "001101100",
3031 => "001101111",
3032 => "001110011",
3033 => "001101001",
3034 => "001100110",
3035 => "001101110",
3036 => "001110000",
3037 => "001100101",
3038 => "001101111",
3039 => "001101011",
3040 => "001101000",
3041 => "001101001",
3042 => "001101010",
3043 => "001101000",
3044 => "001101001",
3045 => "001101100",
3046 => "001101110",
3047 => "001100111",
3048 => "001101011",
3049 => "001100111",
3050 => "001101100",
3051 => "001101010",
3052 => "001101110",
3053 => "001101011",
3054 => "001100111",
3055 => "001101100",
3056 => "001101010",
3057 => "001101011",
3058 => "001101100",
3059 => "001101010",
3060 => "001101000",
3061 => "001100111",
3062 => "001101001",
3063 => "001100110",
3064 => "001100101",
3065 => "001101010",
3066 => "001101010",
3067 => "001101101",
3068 => "001101001",
3069 => "001100110",
3070 => "001101000",
3071 => "001101011",
3072 => "001011101",
3073 => "001100100",
3074 => "001101100",
3075 => "001101001",
3076 => "001110010",
3077 => "001101111",
3078 => "001110010",
3079 => "001110000",
3080 => "001101111",
3081 => "001110010",
3082 => "001110011",
3083 => "001110100",
3084 => "001110010",
3085 => "001110011",
3086 => "001101111",
3087 => "001110111",
3088 => "001110010",
3089 => "001101101",
3090 => "001110000",
3091 => "001101110",
3092 => "001101001",
3093 => "001101011",
3094 => "001101010",
3095 => "001110000",
3096 => "001101110",
3097 => "001101110",
3098 => "001101100",
3099 => "001101100",
3100 => "001101110",
3101 => "001101101",
3102 => "001110001",
3103 => "001110100",
3104 => "001110011",
3105 => "001101100",
3106 => "001101101",
3107 => "001110000",
3108 => "001110010",
3109 => "001110011",
3110 => "001110110",
3111 => "001110100",
3112 => "001110001",
3113 => "001110110",
3114 => "001110001",
3115 => "001101101",
3116 => "001110001",
3117 => "001101111",
3118 => "001101100",
3119 => "001101000",
3120 => "001101001",
3121 => "001101001",
3122 => "001101011",
3123 => "001101110",
3124 => "001101111",
3125 => "001101111",
3126 => "001110001",
3127 => "001101111",
3128 => "001101010",
3129 => "001110001",
3130 => "001110000",
3131 => "001101000",
3132 => "001101011",
3133 => "001101010",
3134 => "001101101",
3135 => "001101100",
3136 => "001101100",
3137 => "001101001",
3138 => "001101001",
3139 => "001101000",
3140 => "001101010",
3141 => "001101001",
3142 => "001100110",
3143 => "001011110",
3144 => "001101011",
3145 => "001101100",
3146 => "001011111",
3147 => "001100010",
3148 => "001101010",
3149 => "001101111",
3150 => "001101011",
3151 => "001101100",
3152 => "001101001",
3153 => "001101011",
3154 => "001101011",
3155 => "001101110",
3156 => "001110011",
3157 => "001110001",
3158 => "001101011",
3159 => "001101011",
3160 => "001101100",
3161 => "001110001",
3162 => "001101011",
3163 => "001101011",
3164 => "001101101",
3165 => "001101100",
3166 => "001100000",
3167 => "001101000",
3168 => "001101111",
3169 => "001101010",
3170 => "001101000",
3171 => "001100101",
3172 => "001110001",
3173 => "001100100",
3174 => "001100110",
3175 => "001101101",
3176 => "001101001",
3177 => "001101001",
3178 => "001101101",
3179 => "001110001",
3180 => "001110011",
3181 => "001101011",
3182 => "001110000",
3183 => "001101110",
3184 => "001100110",
3185 => "001101011",
3186 => "001101001",
3187 => "001100111",
3188 => "001101011",
3189 => "001100110",
3190 => "001100111",
3191 => "001101011",
3192 => "001101010",
3193 => "001101001",
3194 => "001101000",
3195 => "001100110",
3196 => "001100111",
3197 => "001101010",
3198 => "001100110",
3199 => "001100111",
3200 => "001110000",
3201 => "001101110",
3202 => "001101101",
3203 => "001101110",
3204 => "001101111",
3205 => "001110011",
3206 => "001101010",
3207 => "001110010",
3208 => "001101111",
3209 => "001101010",
3210 => "001101100",
3211 => "001100101",
3212 => "001101101",
3213 => "001101101",
3214 => "001101011",
3215 => "001100111",
3216 => "001101011",
3217 => "001101011",
3218 => "001101100",
3219 => "001101101",
3220 => "001101110",
3221 => "001100111",
3222 => "001101001",
3223 => "001100101",
3224 => "001101011",
3225 => "001101000",
3226 => "001101011",
3227 => "001101111",
3228 => "001110001",
3229 => "001110000",
3230 => "001101111",
3231 => "001101110",
3232 => "001101101",
3233 => "001101110",
3234 => "001110000",
3235 => "001110001",
3236 => "001110000",
3237 => "001110001",
3238 => "001110001",
3239 => "001110010",
3240 => "001110001",
3241 => "001110010",
3242 => "001110000",
3243 => "001110000",
3244 => "001110000",
3245 => "001101110",
3246 => "001101111",
3247 => "001101101",
3248 => "001101111",
3249 => "001101110",
3250 => "001101011",
3251 => "001101101",
3252 => "001101101",
3253 => "001110001",
3254 => "001101100",
3255 => "001101111",
3256 => "001101111",
3257 => "001101011",
3258 => "001101110",
3259 => "001101111",
3260 => "001110010",
3261 => "001101100",
3262 => "001101101",
3263 => "001101101",
3264 => "001101101",
3265 => "001101100",
3266 => "001110001",
3267 => "001101100",
3268 => "001101011",
3269 => "001101001",
3270 => "001101110",
3271 => "001100101",
3272 => "001101000",
3273 => "001101010",
3274 => "001101110",
3275 => "001101111",
3276 => "001101110",
3277 => "001101110",
3278 => "001101101",
3279 => "001101101",
3280 => "001101000",
3281 => "001101110",
3282 => "001101111",
3283 => "001101101",
3284 => "001110000",
3285 => "001101111",
3286 => "001101110",
3287 => "001110010",
3288 => "001110001",
3289 => "001101111",
3290 => "001101111",
3291 => "001110001",
3292 => "001110010",
3293 => "001110000",
3294 => "001101110",
3295 => "001110010",
3296 => "001101110",
3297 => "001101111",
3298 => "001110001",
3299 => "001101101",
3300 => "001101011",
3301 => "001110010",
3302 => "001110010",
3303 => "001101010",
3304 => "001110000",
3305 => "001101111",
3306 => "001110010",
3307 => "001101111",
3308 => "001110001",
3309 => "001101110",
3310 => "001101001",
3311 => "001101111",
3312 => "001110001",
3313 => "001101111",
3314 => "001101110",
3315 => "001101110",
3316 => "001101101",
3317 => "001101001",
3318 => "001101110",
3319 => "001101101",
3320 => "001101111",
3321 => "001101111",
3322 => "001110000",
3323 => "001101011",
3324 => "001100110",
3325 => "001101011",
3326 => "001101000",
3327 => "001100100",
3328 => "001110001",
3329 => "001101111",
3330 => "001101110",
3331 => "001101110",
3332 => "001101101",
3333 => "001101011",
3334 => "001101111",
3335 => "001110000",
3336 => "001110010",
3337 => "001101010",
3338 => "001100111",
3339 => "001101000",
3340 => "001101010",
3341 => "001101000",
3342 => "001100111",
3343 => "001100011",
3344 => "001101010",
3345 => "001100111",
3346 => "001101010",
3347 => "001101100",
3348 => "001101010",
3349 => "001101011",
3350 => "001101001",
3351 => "001101101",
3352 => "001101101",
3353 => "001101100",
3354 => "001101101",
3355 => "001101000",
3356 => "001101101",
3357 => "001101100",
3358 => "001101010",
3359 => "001101010",
3360 => "001101100",
3361 => "001101110",
3362 => "001101111",
3363 => "001101001",
3364 => "001101111",
3365 => "001101110",
3366 => "001101110",
3367 => "001101111",
3368 => "001110000",
3369 => "001110011",
3370 => "001110000",
3371 => "001101111",
3372 => "001101110",
3373 => "001110010",
3374 => "001110011",
3375 => "001110010",
3376 => "001101110",
3377 => "001101111",
3378 => "001101101",
3379 => "001110000",
3380 => "001101101",
3381 => "001110000",
3382 => "001101101",
3383 => "001110010",
3384 => "001110000",
3385 => "001110001",
3386 => "001110010",
3387 => "001101111",
3388 => "001101111",
3389 => "001110001",
3390 => "001101101",
3391 => "001101111",
3392 => "001110010",
3393 => "001101111",
3394 => "001110000",
3395 => "001101110",
3396 => "001101110",
3397 => "001101101",
3398 => "001101110",
3399 => "001101110",
3400 => "001101100",
3401 => "001101010",
3402 => "001101111",
3403 => "001101100",
3404 => "001101010",
3405 => "001101110",
3406 => "001101100",
3407 => "001101000",
3408 => "001101001",
3409 => "001100100",
3410 => "001101001",
3411 => "001100100",
3412 => "001101001",
3413 => "001100100",
3414 => "001101011",
3415 => "001101001",
3416 => "001101101",
3417 => "001101001",
3418 => "001101001",
3419 => "001100100",
3420 => "001101011",
3421 => "001101011",
3422 => "001101100",
3423 => "001101011",
3424 => "001101111",
3425 => "001101001",
3426 => "001101010",
3427 => "001101001",
3428 => "001101100",
3429 => "001101101",
3430 => "001100110",
3431 => "001101010",
3432 => "001101111",
3433 => "001101010",
3434 => "001101101",
3435 => "001100111",
3436 => "001101010",
3437 => "001101010",
3438 => "001101011",
3439 => "001100111",
3440 => "001100111",
3441 => "001101001",
3442 => "001100110",
3443 => "001101000",
3444 => "001101000",
3445 => "001101000",
3446 => "001100101",
3447 => "001100101",
3448 => "001100110",
3449 => "001100101",
3450 => "001101000",
3451 => "001101000",
3452 => "001100111",
3453 => "001100100",
3454 => "001100011",
3455 => "001100110",
3456 => "001101101",
3457 => "001101100",
3458 => "001101010",
3459 => "001101011",
3460 => "001100110",
3461 => "001011110",
3462 => "001100111",
3463 => "001100011",
3464 => "001100101",
3465 => "001101001",
3466 => "001100111",
3467 => "001100111",
3468 => "001101000",
3469 => "001100101",
3470 => "001101001",
3471 => "001101000",
3472 => "001101001",
3473 => "001101000",
3474 => "001101100",
3475 => "001101100",
3476 => "001101100",
3477 => "001100111",
3478 => "001101100",
3479 => "001101110",
3480 => "001101100",
3481 => "001101011",
3482 => "001101101",
3483 => "001101111",
3484 => "001110000",
3485 => "001101101",
3486 => "001101111",
3487 => "001101111",
3488 => "001110000",
3489 => "001101100",
3490 => "001101011",
3491 => "001101000",
3492 => "001101011",
3493 => "001101010",
3494 => "001101000",
3495 => "001101011",
3496 => "001101111",
3497 => "001101110",
3498 => "001101110",
3499 => "001101111",
3500 => "001101110",
3501 => "001101010",
3502 => "001101000",
3503 => "001101010",
3504 => "001100111",
3505 => "001100111",
3506 => "001100111",
3507 => "001100101",
3508 => "001101011",
3509 => "001101011",
3510 => "001101010",
3511 => "001101010",
3512 => "001101010",
3513 => "001101101",
3514 => "001101011",
3515 => "001101001",
3516 => "001101100",
3517 => "001101010",
3518 => "001101011",
3519 => "001101001",
3520 => "001101001",
3521 => "001101001",
3522 => "001101010",
3523 => "001101011",
3524 => "001101010",
3525 => "001101011",
3526 => "001100111",
3527 => "001101010",
3528 => "001101001",
3529 => "001101011",
3530 => "001101011",
3531 => "001110010",
3532 => "001101011",
3533 => "001101000",
3534 => "001100111",
3535 => "001101000",
3536 => "001101010",
3537 => "001100101",
3538 => "001100011",
3539 => "001011110",
3540 => "001101001",
3541 => "001100011",
3542 => "001101010",
3543 => "001101100",
3544 => "001100110",
3545 => "001101100",
3546 => "001100111",
3547 => "001101000",
3548 => "001100010",
3549 => "001100011",
3550 => "001100110",
3551 => "001100011",
3552 => "001101011",
3553 => "001100111",
3554 => "001101010",
3555 => "001101000",
3556 => "001100111",
3557 => "001100110",
3558 => "001101001",
3559 => "001100100",
3560 => "001100100",
3561 => "001100101",
3562 => "001100001",
3563 => "001100100",
3564 => "001100100",
3565 => "001100100",
3566 => "001100011",
3567 => "001100101",
3568 => "001100110",
3569 => "001100011",
3570 => "001100101",
3571 => "001100100",
3572 => "001100100",
3573 => "001100011",
3574 => "001100111",
3575 => "001100100",
3576 => "001101011",
3577 => "001100101",
3578 => "001100011",
3579 => "001011101",
3580 => "001100000",
3581 => "001100100",
3582 => "001011111",
3583 => "001100010",
3584 => "001100101",
3585 => "001100001",
3586 => "001100110",
3587 => "001100100",
3588 => "001100100",
3589 => "001101000",
3590 => "001100100",
3591 => "001100100",
3592 => "001100111",
3593 => "001100111",
3594 => "001101100",
3595 => "001101011",
3596 => "001101000",
3597 => "001101000",
3598 => "001101101",
3599 => "001101001",
3600 => "001101011",
3601 => "001101001",
3602 => "001100101",
3603 => "001101010",
3604 => "001101010",
3605 => "001101100",
3606 => "001101111",
3607 => "001101111",
3608 => "001101101",
3609 => "001101101",
3610 => "001101100",
3611 => "001101011",
3612 => "001101101",
3613 => "001101100",
3614 => "001101100",
3615 => "001101101",
3616 => "001101100",
3617 => "001101101",
3618 => "001101001",
3619 => "001101010",
3620 => "001101100",
3621 => "001101101",
3622 => "001101100",
3623 => "001101101",
3624 => "001101111",
3625 => "001110000",
3626 => "001101110",
3627 => "001101011",
3628 => "001101001",
3629 => "001101001",
3630 => "001101000",
3631 => "001101010",
3632 => "001100100",
3633 => "001101001",
3634 => "001101010",
3635 => "001101011",
3636 => "001101110",
3637 => "001101100",
3638 => "001101010",
3639 => "001101101",
3640 => "001110000",
3641 => "001101110",
3642 => "001101110",
3643 => "001101101",
3644 => "001101100",
3645 => "001110001",
3646 => "001101110",
3647 => "001101000",
3648 => "001101100",
3649 => "001101100",
3650 => "001101000",
3651 => "001100111",
3652 => "001100111",
3653 => "001100101",
3654 => "001100110",
3655 => "001101000",
3656 => "001100101",
3657 => "001100011",
3658 => "001101001",
3659 => "001101011",
3660 => "001101011",
3661 => "001100110",
3662 => "001101100",
3663 => "001101001",
3664 => "001100111",
3665 => "001100101",
3666 => "001100110",
3667 => "001101000",
3668 => "001101000",
3669 => "001101011",
3670 => "001100111",
3671 => "001101010",
3672 => "001101000",
3673 => "001101000",
3674 => "001101010",
3675 => "001100110",
3676 => "001100101",
3677 => "001100110",
3678 => "001101001",
3679 => "001100110",
3680 => "001100100",
3681 => "001100110",
3682 => "001100010",
3683 => "001100000",
3684 => "001100101",
3685 => "001100101",
3686 => "001101001",
3687 => "001100101",
3688 => "001100101",
3689 => "001100111",
3690 => "001100110",
3691 => "001100111",
3692 => "001100000",
3693 => "001100110",
3694 => "001100000",
3695 => "001100100",
3696 => "001100001",
3697 => "001100101",
3698 => "001100001",
3699 => "001011110",
3700 => "001100011",
3701 => "001100110",
3702 => "001100010",
3703 => "001100100",
3704 => "001100001",
3705 => "001100010",
3706 => "001100000",
3707 => "001011100",
3708 => "001011110",
3709 => "001011101",
3710 => "001011011",
3711 => "001011101",
3712 => "001101000",
3713 => "001100011",
3714 => "001100001",
3715 => "001100110",
3716 => "001100110",
3717 => "001100101",
3718 => "001100100",
3719 => "001100110",
3720 => "001100100",
3721 => "001100111",
3722 => "001100011",
3723 => "001101000",
3724 => "001100101",
3725 => "001100111",
3726 => "001101011",
3727 => "001101100",
3728 => "001101001",
3729 => "001101000",
3730 => "001101101",
3731 => "001101011",
3732 => "001101101",
3733 => "001101011",
3734 => "001101101",
3735 => "001101100",
3736 => "001101110",
3737 => "001101110",
3738 => "001101011",
3739 => "001101110",
3740 => "001101100",
3741 => "001101111",
3742 => "001101100",
3743 => "001101001",
3744 => "001101101",
3745 => "001101010",
3746 => "001101010",
3747 => "001100111",
3748 => "001100111",
3749 => "001101111",
3750 => "001101100",
3751 => "001101100",
3752 => "001101111",
3753 => "001101111",
3754 => "001101111",
3755 => "001101110",
3756 => "001101100",
3757 => "001101011",
3758 => "001101001",
3759 => "001101001",
3760 => "001101100",
3761 => "001101100",
3762 => "001101100",
3763 => "001101101",
3764 => "001101011",
3765 => "001101100",
3766 => "001101110",
3767 => "001110000",
3768 => "001101110",
3769 => "001101110",
3770 => "001101111",
3771 => "001101100",
3772 => "001101110",
3773 => "001101011",
3774 => "001101111",
3775 => "001101010",
3776 => "001101010",
3777 => "001101011",
3778 => "001101000",
3779 => "001101011",
3780 => "001101010",
3781 => "001101010",
3782 => "001101010",
3783 => "001100111",
3784 => "001101011",
3785 => "001100111",
3786 => "001101001",
3787 => "001100101",
3788 => "001101100",
3789 => "001101011",
3790 => "001101000",
3791 => "001101100",
3792 => "001100111",
3793 => "001101000",
3794 => "001101001",
3795 => "001100011",
3796 => "001101010",
3797 => "001100110",
3798 => "001101000",
3799 => "001100101",
3800 => "001100111",
3801 => "001101100",
3802 => "001101010",
3803 => "001100111",
3804 => "001100101",
3805 => "001100110",
3806 => "001100111",
3807 => "001011110",
3808 => "001100010",
3809 => "001100110",
3810 => "001100111",
3811 => "001100111",
3812 => "001100011",
3813 => "001100011",
3814 => "001100111",
3815 => "001100011",
3816 => "001100101",
3817 => "001100100",
3818 => "001100011",
3819 => "001100000",
3820 => "001100000",
3821 => "001100011",
3822 => "001100010",
3823 => "001011111",
3824 => "001100001",
3825 => "001100000",
3826 => "001100011",
3827 => "001100100",
3828 => "001100110",
3829 => "001100001",
3830 => "001100010",
3831 => "001100011",
3832 => "001100001",
3833 => "001100001",
3834 => "001011110",
3835 => "001100010",
3836 => "001011010",
3837 => "001011101",
3838 => "001011100",
3839 => "001011100",
3840 => "001100101",
3841 => "001100101",
3842 => "001101001",
3843 => "001100110",
3844 => "001100001",
3845 => "001100110",
3846 => "001101001",
3847 => "001100001",
3848 => "001100100",
3849 => "001011111",
3850 => "001100101",
3851 => "001100111",
3852 => "001101010",
3853 => "001100100",
3854 => "001100010",
3855 => "001101000",
3856 => "001101101",
3857 => "001101011",
3858 => "001101011",
3859 => "001101101",
3860 => "001101011",
3861 => "001101011",
3862 => "001100100",
3863 => "001101011",
3864 => "001101011",
3865 => "001100111",
3866 => "001101110",
3867 => "001101011",
3868 => "001101001",
3869 => "001100011",
3870 => "001100010",
3871 => "001101000",
3872 => "001101000",
3873 => "001100110",
3874 => "001101110",
3875 => "001101111",
3876 => "001101100",
3877 => "001101010",
3878 => "001101001",
3879 => "001101011",
3880 => "001101110",
3881 => "001101110",
3882 => "001101010",
3883 => "001101101",
3884 => "001101100",
3885 => "001101110",
3886 => "001101100",
3887 => "001101110",
3888 => "001101100",
3889 => "001101101",
3890 => "001101010",
3891 => "001101010",
3892 => "001101100",
3893 => "001101101",
3894 => "001101101",
3895 => "001101100",
3896 => "001101101",
3897 => "001101111",
3898 => "001110000",
3899 => "001101110",
3900 => "001101100",
3901 => "001101101",
3902 => "001101011",
3903 => "001101011",
3904 => "001101010",
3905 => "001100110",
3906 => "001100101",
3907 => "001101001",
3908 => "001101011",
3909 => "001101011",
3910 => "001100111",
3911 => "001101110",
3912 => "001101110",
3913 => "001100111",
3914 => "001101001",
3915 => "001101100",
3916 => "001101010",
3917 => "001101111",
3918 => "001101000",
3919 => "001100110",
3920 => "001101011",
3921 => "001101100",
3922 => "001100100",
3923 => "001100111",
3924 => "001101000",
3925 => "001100101",
3926 => "001100110",
3927 => "001101011",
3928 => "001101010",
3929 => "001100111",
3930 => "001100110",
3931 => "001100111",
3932 => "001100010",
3933 => "001100111",
3934 => "001100111",
3935 => "001101011",
3936 => "001101011",
3937 => "001100110",
3938 => "001101000",
3939 => "001100110",
3940 => "001100100",
3941 => "001100101",
3942 => "001011110",
3943 => "001100011",
3944 => "001100011",
3945 => "001100101",
3946 => "001100011",
3947 => "001100100",
3948 => "001100011",
3949 => "001100001",
3950 => "001100100",
3951 => "001100010",
3952 => "001100001",
3953 => "001100001",
3954 => "001100001",
3955 => "001100010",
3956 => "001100100",
3957 => "001100001",
3958 => "001100000",
3959 => "001100010",
3960 => "001011110",
3961 => "001011101",
3962 => "001011111",
3963 => "001100101",
3964 => "001011111",
3965 => "001100001",
3966 => "001011111",
3967 => "001011100",
3968 => "001011111",
3969 => "001100101",
3970 => "001100010",
3971 => "001100011",
3972 => "001100010",
3973 => "001011111",
3974 => "001100001",
3975 => "001100001",
3976 => "001100000",
3977 => "001100010",
3978 => "001011111",
3979 => "001011010",
3980 => "001101000",
3981 => "001101001",
3982 => "001100110",
3983 => "001100001",
3984 => "001100011",
3985 => "001101000",
3986 => "001100111",
3987 => "001100111",
3988 => "001100111",
3989 => "001101011",
3990 => "001101010",
3991 => "001101010",
3992 => "001101001",
3993 => "001101001",
3994 => "001101001",
3995 => "001101011",
3996 => "001101110",
3997 => "001101010",
3998 => "001100100",
3999 => "001101011",
4000 => "001101100",
4001 => "001101100",
4002 => "001101010",
4003 => "001101101",
4004 => "001101100",
4005 => "001101011",
4006 => "001101000",
4007 => "001101010",
4008 => "001101101",
4009 => "001101101",
4010 => "001101010",
4011 => "001101001",
4012 => "001101001",
4013 => "001100101",
4014 => "001101010",
4015 => "001100111",
4016 => "001101000",
4017 => "001100111",
4018 => "001110001",
4019 => "001100100",
4020 => "001101001",
4021 => "001100111",
4022 => "001101011",
4023 => "001101101",
4024 => "001101001",
4025 => "001101010",
4026 => "001101001",
4027 => "001101001",
4028 => "001101000",
4029 => "001100101",
4030 => "001100101",
4031 => "001100101",
4032 => "001101000",
4033 => "001101001",
4034 => "001100111",
4035 => "001101011",
4036 => "001101011",
4037 => "001101001",
4038 => "001101011",
4039 => "001101011",
4040 => "001101100",
4041 => "001101100",
4042 => "001101000",
4043 => "001100111",
4044 => "001101000",
4045 => "001101000",
4046 => "001101000",
4047 => "001101010",
4048 => "001100100",
4049 => "001101001",
4050 => "001100111",
4051 => "001101000",
4052 => "001011111",
4053 => "001101010",
4054 => "001100110",
4055 => "001100101",
4056 => "001100100",
4057 => "001101000",
4058 => "001100110",
4059 => "001100100",
4060 => "001100110",
4061 => "001101001",
4062 => "001101110",
4063 => "001100111",
4064 => "001100110",
4065 => "001101001",
4066 => "001100110",
4067 => "001101001",
4068 => "001100110",
4069 => "001100001",
4070 => "001100110",
4071 => "001100100",
4072 => "001100100",
4073 => "001100100",
4074 => "001100100",
4075 => "001100110",
4076 => "001100101",
4077 => "001100110",
4078 => "001100110",
4079 => "001100111",
4080 => "001100111",
4081 => "001100101",
4082 => "001100100",
4083 => "001100101",
4084 => "001100010",
4085 => "001100001",
4086 => "001100010",
4087 => "001011111",
4088 => "001011111",
4089 => "001011101",
4090 => "001011101",
4091 => "001011111",
4092 => "001100000",
4093 => "001011111",
4094 => "001100000",
4095 => "001011010",
4096 => "001011111",
4097 => "001011110",
4098 => "001100001",
4099 => "001100100",
4100 => "001100000",
4101 => "001100011",
4102 => "001100101",
4103 => "001100101",
4104 => "001100111",
4105 => "001100010",
4106 => "001101000",
4107 => "001100111",
4108 => "001101010",
4109 => "001101100",
4110 => "001101010",
4111 => "001101101",
4112 => "001101011",
4113 => "001101001",
4114 => "001101100",
4115 => "001100110",
4116 => "001101000",
4117 => "001100111",
4118 => "001100101",
4119 => "001101100",
4120 => "001100111",
4121 => "001101000",
4122 => "001100101",
4123 => "001011111",
4124 => "001100111",
4125 => "001100110",
4126 => "001101111",
4127 => "001101011",
4128 => "001101000",
4129 => "001101001",
4130 => "001101001",
4131 => "001100001",
4132 => "001101101",
4133 => "001100101",
4134 => "001100101",
4135 => "001101001",
4136 => "001101001",
4137 => "001100101",
4138 => "001100110",
4139 => "001011111",
4140 => "001100110",
4141 => "001100101",
4142 => "001100110",
4143 => "001100100",
4144 => "001100101",
4145 => "001110100",
4146 => "010000001",
4147 => "001101000",
4148 => "001101000",
4149 => "001101000",
4150 => "001100100",
4151 => "001101000",
4152 => "001100101",
4153 => "001100110",
4154 => "001100010",
4155 => "001101011",
4156 => "001101011",
4157 => "001101101",
4158 => "001101010",
4159 => "001101001",
4160 => "001100111",
4161 => "001101000",
4162 => "001100111",
4163 => "001101011",
4164 => "001101111",
4165 => "001101010",
4166 => "001101011",
4167 => "001101010",
4168 => "001101011",
4169 => "001101011",
4170 => "001101110",
4171 => "001101110",
4172 => "001101000",
4173 => "001101001",
4174 => "001101010",
4175 => "001100110",
4176 => "001100111",
4177 => "001100100",
4178 => "001100110",
4179 => "001100110",
4180 => "001100110",
4181 => "001100110",
4182 => "001100100",
4183 => "001100110",
4184 => "001101001",
4185 => "001101100",
4186 => "001101100",
4187 => "001100110",
4188 => "001100011",
4189 => "001101001",
4190 => "001101010",
4191 => "001101011",
4192 => "001101011",
4193 => "001101010",
4194 => "001100111",
4195 => "001100010",
4196 => "001100101",
4197 => "001100111",
4198 => "001101010",
4199 => "001100111",
4200 => "001100011",
4201 => "001101000",
4202 => "001100101",
4203 => "001100001",
4204 => "001011011",
4205 => "001100100",
4206 => "001100000",
4207 => "001100001",
4208 => "001100010",
4209 => "001100010",
4210 => "001011110",
4211 => "001011100",
4212 => "001100010",
4213 => "001100001",
4214 => "001100001",
4215 => "001100001",
4216 => "001011111",
4217 => "001100000",
4218 => "001100000",
4219 => "001100011",
4220 => "001100010",
4221 => "001011011",
4222 => "001011100",
4223 => "001100001",
4224 => "001100100",
4225 => "001100010",
4226 => "001100101",
4227 => "001100000",
4228 => "001100001",
4229 => "001100011",
4230 => "001100010",
4231 => "001100101",
4232 => "001011111",
4233 => "001101001",
4234 => "001100111",
4235 => "001101000",
4236 => "001100111",
4237 => "001100100",
4238 => "001100111",
4239 => "001101010",
4240 => "001101000",
4241 => "001101001",
4242 => "001101000",
4243 => "001101000",
4244 => "001100101",
4245 => "001100110",
4246 => "001100100",
4247 => "001011111",
4248 => "001100010",
4249 => "001101010",
4250 => "001100011",
4251 => "001100101",
4252 => "001101001",
4253 => "001101011",
4254 => "001101010",
4255 => "001100100",
4256 => "001100001",
4257 => "001011111",
4258 => "001100011",
4259 => "001100101",
4260 => "001100101",
4261 => "001100111",
4262 => "001100011",
4263 => "001101001",
4264 => "001101011",
4265 => "001101010",
4266 => "001100110",
4267 => "001101011",
4268 => "001100101",
4269 => "001101000",
4270 => "001100110",
4271 => "001101010",
4272 => "001110001",
4273 => "010100110",
4274 => "010110000",
4275 => "010001111",
4276 => "001011101",
4277 => "001100001",
4278 => "001100110",
4279 => "001101000",
4280 => "001100111",
4281 => "001100111",
4282 => "001101010",
4283 => "001101111",
4284 => "001101011",
4285 => "001101111",
4286 => "001101001",
4287 => "001101011",
4288 => "001100110",
4289 => "001101101",
4290 => "001101010",
4291 => "001101101",
4292 => "001101110",
4293 => "001101110",
4294 => "001101111",
4295 => "001101101",
4296 => "001101011",
4297 => "001101011",
4298 => "001101100",
4299 => "001101100",
4300 => "001101100",
4301 => "001101011",
4302 => "001101101",
4303 => "001101001",
4304 => "001101011",
4305 => "001101010",
4306 => "001101100",
4307 => "001100111",
4308 => "001100111",
4309 => "001101001",
4310 => "001101010",
4311 => "001100110",
4312 => "001101011",
4313 => "001101110",
4314 => "001101100",
4315 => "001100100",
4316 => "001101010",
4317 => "001101100",
4318 => "001101000",
4319 => "001100101",
4320 => "001100010",
4321 => "001100101",
4322 => "001100110",
4323 => "001100110",
4324 => "001100010",
4325 => "001100101",
4326 => "001100010",
4327 => "001100010",
4328 => "001100011",
4329 => "001100001",
4330 => "001100001",
4331 => "001011111",
4332 => "001100011",
4333 => "001100010",
4334 => "001011100",
4335 => "001011101",
4336 => "001011111",
4337 => "001101000",
4338 => "001100000",
4339 => "001100000",
4340 => "001100100",
4341 => "001100100",
4342 => "001101000",
4343 => "001100001",
4344 => "001011110",
4345 => "001100010",
4346 => "001100101",
4347 => "001101001",
4348 => "001100011",
4349 => "001011110",
4350 => "001011100",
4351 => "001011010",
4352 => "001011111",
4353 => "001011101",
4354 => "001100011",
4355 => "001011111",
4356 => "001100101",
4357 => "001100101",
4358 => "001100110",
4359 => "001100101",
4360 => "001101010",
4361 => "001100101",
4362 => "001101001",
4363 => "001100100",
4364 => "001101101",
4365 => "001101000",
4366 => "001100110",
4367 => "001101101",
4368 => "001101100",
4369 => "001101011",
4370 => "001100110",
4371 => "001100101",
4372 => "001101001",
4373 => "001100110",
4374 => "001100100",
4375 => "001101001",
4376 => "001100100",
4377 => "001100101",
4378 => "001011111",
4379 => "001101000",
4380 => "001101001",
4381 => "001101000",
4382 => "001100001",
4383 => "001101000",
4384 => "001100100",
4385 => "001100111",
4386 => "001101001",
4387 => "001100010",
4388 => "001100001",
4389 => "001100010",
4390 => "001011100",
4391 => "001101001",
4392 => "001101010",
4393 => "001101011",
4394 => "001101101",
4395 => "001101110",
4396 => "001101000",
4397 => "001101100",
4398 => "001101111",
4399 => "001101011",
4400 => "010011101",
4401 => "011001010",
4402 => "010000000",
4403 => "001100000",
4404 => "001101111",
4405 => "001110001",
4406 => "001110010",
4407 => "001101010",
4408 => "001101100",
4409 => "001101000",
4410 => "001100111",
4411 => "001100011",
4412 => "001101011",
4413 => "001100111",
4414 => "001101010",
4415 => "001100110",
4416 => "001101001",
4417 => "001101011",
4418 => "001101100",
4419 => "001100101",
4420 => "001100110",
4421 => "001101010",
4422 => "001101001",
4423 => "001101010",
4424 => "001101110",
4425 => "001110000",
4426 => "001101001",
4427 => "001101000",
4428 => "001101010",
4429 => "001101110",
4430 => "001100100",
4431 => "001101011",
4432 => "001101111",
4433 => "001101100",
4434 => "001101110",
4435 => "001101100",
4436 => "001101100",
4437 => "001100111",
4438 => "001101000",
4439 => "001101010",
4440 => "001101101",
4441 => "010000010",
4442 => "010011010",
4443 => "011000010",
4444 => "001101001",
4445 => "001101100",
4446 => "001101100",
4447 => "001101010",
4448 => "001100110",
4449 => "001101000",
4450 => "001100110",
4451 => "001100100",
4452 => "001100100",
4453 => "001100001",
4454 => "001100101",
4455 => "001100101",
4456 => "001100011",
4457 => "001100010",
4458 => "001100010",
4459 => "001100001",
4460 => "001100001",
4461 => "001100101",
4462 => "001100111",
4463 => "001100100",
4464 => "001101000",
4465 => "001100101",
4466 => "001100010",
4467 => "001100100",
4468 => "001100001",
4469 => "001100001",
4470 => "001100011",
4471 => "001100011",
4472 => "001100011",
4473 => "001100001",
4474 => "001011000",
4475 => "001011110",
4476 => "001011101",
4477 => "001011111",
4478 => "001011111",
4479 => "001011011",
4480 => "001100000",
4481 => "001100100",
4482 => "001100001",
4483 => "001100000",
4484 => "001100000",
4485 => "001100011",
4486 => "001011010",
4487 => "001100100",
4488 => "001100100",
4489 => "001100011",
4490 => "001101010",
4491 => "001100010",
4492 => "001100110",
4493 => "001101010",
4494 => "001101010",
4495 => "001101010",
4496 => "001101000",
4497 => "001101000",
4498 => "001100111",
4499 => "001100101",
4500 => "001100101",
4501 => "001100101",
4502 => "001100110",
4503 => "001100100",
4504 => "001101000",
4505 => "001100110",
4506 => "001100010",
4507 => "001100111",
4508 => "001101000",
4509 => "001100100",
4510 => "001100111",
4511 => "001101000",
4512 => "001101100",
4513 => "001101000",
4514 => "001101100",
4515 => "001101101",
4516 => "001101001",
4517 => "001101000",
4518 => "001101001",
4519 => "001101100",
4520 => "001101010",
4521 => "001101101",
4522 => "001101101",
4523 => "001101111",
4524 => "001101100",
4525 => "001101100",
4526 => "001101110",
4527 => "010101101",
4528 => "011000100",
4529 => "010101111",
4530 => "001011110",
4531 => "001010110",
4532 => "001011011",
4533 => "001100100",
4534 => "001011111",
4535 => "001011010",
4536 => "001101001",
4537 => "001110001",
4538 => "001110000",
4539 => "001101110",
4540 => "001101001",
4541 => "001101011",
4542 => "001101001",
4543 => "001100000",
4544 => "001101010",
4545 => "001101001",
4546 => "001100110",
4547 => "001101011",
4548 => "001101000",
4549 => "001101000",
4550 => "001101010",
4551 => "001101100",
4552 => "001100011",
4553 => "001100101",
4554 => "001101000",
4555 => "001101000",
4556 => "001101011",
4557 => "001101001",
4558 => "001101010",
4559 => "001101010",
4560 => "001100011",
4561 => "001101001",
4562 => "001101010",
4563 => "001101001",
4564 => "001101010",
4565 => "001100111",
4566 => "001101001",
4567 => "001101010",
4568 => "001101101",
4569 => "010010101",
4570 => "010111100",
4571 => "011001111",
4572 => "011011100",
4573 => "001101100",
4574 => "001100110",
4575 => "001100100",
4576 => "001100100",
4577 => "001100001",
4578 => "001100110",
4579 => "001100100",
4580 => "001100100",
4581 => "001100001",
4582 => "001100001",
4583 => "001100010",
4584 => "001011110",
4585 => "001011110",
4586 => "001100101",
4587 => "001100100",
4588 => "001100010",
4589 => "001100010",
4590 => "001100001",
4591 => "001100100",
4592 => "001100000",
4593 => "001011101",
4594 => "001011110",
4595 => "001100001",
4596 => "001100010",
4597 => "001100001",
4598 => "001011110",
4599 => "001011101",
4600 => "001100011",
4601 => "001100010",
4602 => "001100010",
4603 => "001011110",
4604 => "001100001",
4605 => "001010110",
4606 => "001010100",
4607 => "001011011",
4608 => "001100000",
4609 => "001100011",
4610 => "001100001",
4611 => "001100000",
4612 => "001100010",
4613 => "001100100",
4614 => "001100011",
4615 => "001100100",
4616 => "001100110",
4617 => "001101011",
4618 => "001101001",
4619 => "001100011",
4620 => "001100010",
4621 => "001101011",
4622 => "001101011",
4623 => "001101000",
4624 => "001100101",
4625 => "001100111",
4626 => "001101010",
4627 => "001100111",
4628 => "001101010",
4629 => "001101000",
4630 => "001101001",
4631 => "001100101",
4632 => "001100111",
4633 => "001100111",
4634 => "001101010",
4635 => "001101010",
4636 => "001101100",
4637 => "001101001",
4638 => "001101101",
4639 => "001101101",
4640 => "001101011",
4641 => "001101001",
4642 => "001101001",
4643 => "001101011",
4644 => "001101010",
4645 => "001101000",
4646 => "001101100",
4647 => "001101101",
4648 => "001101011",
4649 => "001101001",
4650 => "001101111",
4651 => "001101110",
4652 => "001100111",
4653 => "001101100",
4654 => "010011111",
4655 => "011010100",
4656 => "011001011",
4657 => "001101010",
4658 => "001100100",
4659 => "001100111",
4660 => "001100110",
4661 => "001100010",
4662 => "001011000",
4663 => "001011010",
4664 => "001011100",
4665 => "001100100",
4666 => "001011000",
4667 => "001011001",
4668 => "001001010",
4669 => "001101010",
4670 => "001110000",
4671 => "001101111",
4672 => "001100111",
4673 => "001100101",
4674 => "001100101",
4675 => "001101001",
4676 => "001101010",
4677 => "001101101",
4678 => "001101101",
4679 => "001101110",
4680 => "001101001",
4681 => "001101001",
4682 => "001101101",
4683 => "001101001",
4684 => "001100100",
4685 => "001101000",
4686 => "001101001",
4687 => "001100101",
4688 => "001100111",
4689 => "001101100",
4690 => "001101000",
4691 => "001100101",
4692 => "001100101",
4693 => "001100010",
4694 => "001101010",
4695 => "001100101",
4696 => "010000001",
4697 => "010100000",
4698 => "011101111",
4699 => "010101111",
4700 => "011101011",
4701 => "010011101",
4702 => "001100100",
4703 => "001100010",
4704 => "001100110",
4705 => "001100111",
4706 => "001100011",
4707 => "001100100",
4708 => "001101010",
4709 => "001100111",
4710 => "001100100",
4711 => "001100000",
4712 => "001100001",
4713 => "001100100",
4714 => "001100110",
4715 => "001100110",
4716 => "001100110",
4717 => "001100100",
4718 => "001100111",
4719 => "001101000",
4720 => "001100110",
4721 => "001100101",
4722 => "001100010",
4723 => "001100001",
4724 => "001100001",
4725 => "001011110",
4726 => "001100001",
4727 => "001011100",
4728 => "001010111",
4729 => "001011001",
4730 => "001011100",
4731 => "001011011",
4732 => "001011001",
4733 => "001011110",
4734 => "001011001",
4735 => "001011001",
4736 => "001011110",
4737 => "001011110",
4738 => "001100011",
4739 => "001100011",
4740 => "001100001",
4741 => "001100001",
4742 => "001100111",
4743 => "001011111",
4744 => "001100101",
4745 => "001100100",
4746 => "001100100",
4747 => "001100110",
4748 => "001100101",
4749 => "001101011",
4750 => "001101000",
4751 => "001100100",
4752 => "001101011",
4753 => "001100101",
4754 => "001100100",
4755 => "001101011",
4756 => "001101011",
4757 => "001101111",
4758 => "001101111",
4759 => "001101100",
4760 => "001101001",
4761 => "001101010",
4762 => "001101100",
4763 => "001101011",
4764 => "001101010",
4765 => "001101011",
4766 => "001101101",
4767 => "001101011",
4768 => "001101110",
4769 => "001101110",
4770 => "001101111",
4771 => "001110001",
4772 => "001110010",
4773 => "001101111",
4774 => "001110001",
4775 => "001101101",
4776 => "001101101",
4777 => "001101110",
4778 => "001101111",
4779 => "001101111",
4780 => "001110001",
4781 => "010000001",
4782 => "011010101",
4783 => "011001100",
4784 => "001111011",
4785 => "001100110",
4786 => "001100101",
4787 => "001100100",
4788 => "001100010",
4789 => "001100010",
4790 => "001100101",
4791 => "001100100",
4792 => "001011110",
4793 => "001011001",
4794 => "001011011",
4795 => "001100000",
4796 => "001100100",
4797 => "001011100",
4798 => "001011110",
4799 => "001011101",
4800 => "001011100",
4801 => "001100010",
4802 => "001011111",
4803 => "001101011",
4804 => "001101010",
4805 => "001101010",
4806 => "001100111",
4807 => "001100100",
4808 => "001100101",
4809 => "001100011",
4810 => "001100101",
4811 => "001100100",
4812 => "001100111",
4813 => "001100111",
4814 => "001101001",
4815 => "001100111",
4816 => "001100101",
4817 => "001100110",
4818 => "001100100",
4819 => "001100010",
4820 => "001100100",
4821 => "001100100",
4822 => "001101000",
4823 => "001110111",
4824 => "010000100",
4825 => "010111000",
4826 => "011010011",
4827 => "001111001",
4828 => "011101111",
4829 => "011100110",
4830 => "001101110",
4831 => "001100111",
4832 => "001100011",
4833 => "001100100",
4834 => "001100111",
4835 => "001100101",
4836 => "001100000",
4837 => "001100011",
4838 => "001100011",
4839 => "001100011",
4840 => "001100011",
4841 => "001100101",
4842 => "001100011",
4843 => "001100101",
4844 => "001100110",
4845 => "001100001",
4846 => "001011110",
4847 => "001100001",
4848 => "001011100",
4849 => "001011101",
4850 => "001100010",
4851 => "001100000",
4852 => "001100001",
4853 => "001011011",
4854 => "001011100",
4855 => "001011101",
4856 => "001011101",
4857 => "001011101",
4858 => "001100100",
4859 => "001011101",
4860 => "001011110",
4861 => "001011111",
4862 => "001011101",
4863 => "001011111",
4864 => "001100011",
4865 => "001100001",
4866 => "001100000",
4867 => "001100001",
4868 => "001100100",
4869 => "001100010",
4870 => "001011100",
4871 => "001100010",
4872 => "001100010",
4873 => "001100000",
4874 => "001100100",
4875 => "001100100",
4876 => "001101000",
4877 => "001100010",
4878 => "001100010",
4879 => "001100101",
4880 => "001100110",
4881 => "001100100",
4882 => "001100010",
4883 => "001101000",
4884 => "001101101",
4885 => "001101001",
4886 => "001101011",
4887 => "001101011",
4888 => "001101101",
4889 => "001101011",
4890 => "001101010",
4891 => "001101001",
4892 => "001101011",
4893 => "001101110",
4894 => "001110000",
4895 => "001101101",
4896 => "001101111",
4897 => "001101100",
4898 => "001101100",
4899 => "001101100",
4900 => "001101010",
4901 => "001101010",
4902 => "001101000",
4903 => "001101011",
4904 => "001101111",
4905 => "001101010",
4906 => "001101100",
4907 => "001101110",
4908 => "001101001",
4909 => "011001100",
4910 => "011011000",
4911 => "010000001",
4912 => "001100101",
4913 => "001100100",
4914 => "001100011",
4915 => "001100010",
4916 => "001100100",
4917 => "001100010",
4918 => "001100011",
4919 => "001100101",
4920 => "001100101",
4921 => "001100010",
4922 => "001100010",
4923 => "001011100",
4924 => "001011101",
4925 => "001011100",
4926 => "001011000",
4927 => "001011011",
4928 => "001011011",
4929 => "001011000",
4930 => "001011011",
4931 => "001011011",
4932 => "001011101",
4933 => "001011001",
4934 => "001100000",
4935 => "001100010",
4936 => "001101010",
4937 => "001110011",
4938 => "001101010",
4939 => "001101000",
4940 => "001100100",
4941 => "001100010",
4942 => "001100011",
4943 => "001100001",
4944 => "001100010",
4945 => "001100100",
4946 => "001100111",
4947 => "001101000",
4948 => "001100100",
4949 => "001100110",
4950 => "001100110",
4951 => "010011100",
4952 => "010110000",
4953 => "011101000",
4954 => "010111101",
4955 => "001100101",
4956 => "011100110",
4957 => "011100111",
4958 => "001111001",
4959 => "001100111",
4960 => "001100011",
4961 => "001101000",
4962 => "001100010",
4963 => "001100001",
4964 => "001101000",
4965 => "001100110",
4966 => "001011110",
4967 => "001011100",
4968 => "001011110",
4969 => "001011101",
4970 => "001011111",
4971 => "001011111",
4972 => "001011111",
4973 => "001011110",
4974 => "001011111",
4975 => "001011010",
4976 => "001100000",
4977 => "001100001",
4978 => "001100000",
4979 => "001100100",
4980 => "001100011",
4981 => "001100011",
4982 => "001011100",
4983 => "001011010",
4984 => "001011011",
4985 => "001011111",
4986 => "001100000",
4987 => "001100011",
4988 => "001100011",
4989 => "001100010",
4990 => "001100000",
4991 => "001011010",
4992 => "001100100",
4993 => "001100110",
4994 => "001100011",
4995 => "001100011",
4996 => "001100110",
4997 => "001100101",
4998 => "001100110",
4999 => "001100101",
5000 => "001100011",
5001 => "001100110",
5002 => "001101011",
5003 => "001100111",
5004 => "001100101",
5005 => "001101000",
5006 => "001100101",
5007 => "001100110",
5008 => "001101000",
5009 => "001101011",
5010 => "001101101",
5011 => "001101010",
5012 => "001101011",
5013 => "001101010",
5014 => "001100110",
5015 => "001101000",
5016 => "001101010",
5017 => "001101001",
5018 => "001100111",
5019 => "001101000",
5020 => "001100111",
5021 => "001101001",
5022 => "001100111",
5023 => "001101000",
5024 => "001101011",
5025 => "001101001",
5026 => "001101010",
5027 => "001101000",
5028 => "001100011",
5029 => "001100010",
5030 => "001100101",
5031 => "001100101",
5032 => "001100101",
5033 => "001101001",
5034 => "001101001",
5035 => "001101011",
5036 => "010110110",
5037 => "011010010",
5038 => "010010101",
5039 => "001101000",
5040 => "001100111",
5041 => "001100111",
5042 => "001100001",
5043 => "001100011",
5044 => "001100100",
5045 => "001100001",
5046 => "001100010",
5047 => "001100000",
5048 => "001100010",
5049 => "001100010",
5050 => "001100110",
5051 => "001100101",
5052 => "001100001",
5053 => "001100000",
5054 => "001100011",
5055 => "001100011",
5056 => "001100100",
5057 => "001100101",
5058 => "001100000",
5059 => "001010101",
5060 => "001011001",
5061 => "001011001",
5062 => "001010111",
5063 => "001010110",
5064 => "001010111",
5065 => "001011101",
5066 => "001100001",
5067 => "001100100",
5068 => "001101100",
5069 => "001101011",
5070 => "001101011",
5071 => "001101100",
5072 => "001101001",
5073 => "001100110",
5074 => "001100110",
5075 => "001100100",
5076 => "001101000",
5077 => "001101011",
5078 => "001101000",
5079 => "010101110",
5080 => "011000101",
5081 => "011100100",
5082 => "001101111",
5083 => "010101010",
5084 => "011100001",
5085 => "011101000",
5086 => "010001110",
5087 => "001011110",
5088 => "001011111",
5089 => "001011011",
5090 => "001011110",
5091 => "001011111",
5092 => "001011111",
5093 => "001100001",
5094 => "001011111",
5095 => "001011111",
5096 => "001100010",
5097 => "001100001",
5098 => "001011101",
5099 => "001011001",
5100 => "001011100",
5101 => "001011110",
5102 => "001011110",
5103 => "001011100",
5104 => "001011101",
5105 => "001010110",
5106 => "001011100",
5107 => "001100000",
5108 => "001100001",
5109 => "001100001",
5110 => "001100000",
5111 => "001011111",
5112 => "001011111",
5113 => "001011101",
5114 => "001011010",
5115 => "001011110",
5116 => "001100000",
5117 => "001011101",
5118 => "001011111",
5119 => "001011010",
5120 => "001100100",
5121 => "001100100",
5122 => "001100010",
5123 => "001100001",
5124 => "001100010",
5125 => "001011110",
5126 => "001011111",
5127 => "001100101",
5128 => "001100011",
5129 => "001100111",
5130 => "001100100",
5131 => "001101000",
5132 => "001101000",
5133 => "001100111",
5134 => "001100110",
5135 => "001101001",
5136 => "001100101",
5137 => "001100001",
5138 => "001101000",
5139 => "001101001",
5140 => "001101101",
5141 => "001101110",
5142 => "001101010",
5143 => "001101001",
5144 => "001101100",
5145 => "001101100",
5146 => "001101010",
5147 => "001101010",
5148 => "001101010",
5149 => "001101010",
5150 => "001100110",
5151 => "001100111",
5152 => "001101000",
5153 => "001101001",
5154 => "001101100",
5155 => "001101101",
5156 => "001101100",
5157 => "001101101",
5158 => "001101101",
5159 => "001101110",
5160 => "001110001",
5161 => "001101101",
5162 => "001101011",
5163 => "010011100",
5164 => "011010111",
5165 => "010101111",
5166 => "001101010",
5167 => "001100111",
5168 => "001101001",
5169 => "001100011",
5170 => "001100100",
5171 => "001100101",
5172 => "001100011",
5173 => "001100011",
5174 => "001100001",
5175 => "001100011",
5176 => "001100010",
5177 => "001100011",
5178 => "001100011",
5179 => "001011111",
5180 => "001011111",
5181 => "001100001",
5182 => "001100010",
5183 => "001100000",
5184 => "001100100",
5185 => "001100010",
5186 => "001011111",
5187 => "001100010",
5188 => "001100000",
5189 => "001011111",
5190 => "001100010",
5191 => "001100100",
5192 => "001011100",
5193 => "001010110",
5194 => "001011000",
5195 => "001100000",
5196 => "001011000",
5197 => "001011000",
5198 => "001011010",
5199 => "001011010",
5200 => "001100100",
5201 => "001100001",
5202 => "001100101",
5203 => "001100111",
5204 => "001101010",
5205 => "001101001",
5206 => "001110110",
5207 => "010110000",
5208 => "011010111",
5209 => "011101000",
5210 => "001110010",
5211 => "011000001",
5212 => "011101000",
5213 => "011110011",
5214 => "010001011",
5215 => "001101100",
5216 => "001101011",
5217 => "001101000",
5218 => "001101010",
5219 => "001101000",
5220 => "001100110",
5221 => "001100011",
5222 => "001100011",
5223 => "001011110",
5224 => "001100000",
5225 => "001011110",
5226 => "001100010",
5227 => "001100011",
5228 => "001100011",
5229 => "001100001",
5230 => "001100101",
5231 => "001100101",
5232 => "001100101",
5233 => "001100100",
5234 => "001100001",
5235 => "001100001",
5236 => "001100011",
5237 => "001100000",
5238 => "001100010",
5239 => "001100100",
5240 => "001100100",
5241 => "001100011",
5242 => "001100000",
5243 => "001100010",
5244 => "001100000",
5245 => "001100100",
5246 => "001100011",
5247 => "001100100",
5248 => "001100011",
5249 => "001100100",
5250 => "001100110",
5251 => "001100011",
5252 => "001100110",
5253 => "001101100",
5254 => "001100101",
5255 => "001100111",
5256 => "001100110",
5257 => "001101001",
5258 => "001101011",
5259 => "001101001",
5260 => "001100100",
5261 => "001100110",
5262 => "001100110",
5263 => "001100101",
5264 => "001101000",
5265 => "001100110",
5266 => "001101011",
5267 => "001100011",
5268 => "001100010",
5269 => "001100100",
5270 => "001100101",
5271 => "001100010",
5272 => "001100101",
5273 => "001101011",
5274 => "001101000",
5275 => "001100110",
5276 => "001100111",
5277 => "001101001",
5278 => "001101010",
5279 => "001101100",
5280 => "001101101",
5281 => "001101101",
5282 => "001101100",
5283 => "001101101",
5284 => "001101110",
5285 => "001101101",
5286 => "001101100",
5287 => "001101100",
5288 => "001101011",
5289 => "001101010",
5290 => "001111111",
5291 => "011011111",
5292 => "011000111",
5293 => "001101101",
5294 => "001100101",
5295 => "001100110",
5296 => "001100101",
5297 => "001100001",
5298 => "001100010",
5299 => "001100010",
5300 => "001100101",
5301 => "001100001",
5302 => "001100100",
5303 => "001100011",
5304 => "001100011",
5305 => "001100100",
5306 => "001100000",
5307 => "001100001",
5308 => "001100100",
5309 => "001100001",
5310 => "001100001",
5311 => "001100010",
5312 => "001100001",
5313 => "001100000",
5314 => "001100011",
5315 => "001100010",
5316 => "001100001",
5317 => "001100001",
5318 => "001100001",
5319 => "001011111",
5320 => "001100010",
5321 => "001100011",
5322 => "001100110",
5323 => "001100001",
5324 => "001100001",
5325 => "001011101",
5326 => "001010010",
5327 => "001010100",
5328 => "001010101",
5329 => "001010110",
5330 => "001010011",
5331 => "001001110",
5332 => "001000011",
5333 => "001001011",
5334 => "001110101",
5335 => "010110111",
5336 => "011011010",
5337 => "011101101",
5338 => "011101000",
5339 => "011011010",
5340 => "011011111",
5341 => "011100110",
5342 => "001111110",
5343 => "001100111",
5344 => "001100100",
5345 => "001100111",
5346 => "001100111",
5347 => "001100000",
5348 => "001100011",
5349 => "001100110",
5350 => "001100110",
5351 => "001100001",
5352 => "001100011",
5353 => "001100001",
5354 => "001100101",
5355 => "001100001",
5356 => "001011110",
5357 => "001100101",
5358 => "001100010",
5359 => "001011111",
5360 => "001100001",
5361 => "001100010",
5362 => "001100010",
5363 => "001011011",
5364 => "001100001",
5365 => "001100100",
5366 => "001100010",
5367 => "001100101",
5368 => "001100000",
5369 => "001011011",
5370 => "001011100",
5371 => "001011011",
5372 => "001100001",
5373 => "001100000",
5374 => "001011111",
5375 => "001011111",
5376 => "001100000",
5377 => "001100011",
5378 => "001011101",
5379 => "001011011",
5380 => "001100001",
5381 => "001100001",
5382 => "001100001",
5383 => "001011110",
5384 => "001011111",
5385 => "001100001",
5386 => "001100001",
5387 => "001100001",
5388 => "001100010",
5389 => "001100110",
5390 => "001100111",
5391 => "001100111",
5392 => "001100000",
5393 => "001100110",
5394 => "001100101",
5395 => "001100110",
5396 => "001100111",
5397 => "001100101",
5398 => "001101001",
5399 => "001100000",
5400 => "001100101",
5401 => "001100100",
5402 => "001100010",
5403 => "001100001",
5404 => "001100001",
5405 => "001011010",
5406 => "001100101",
5407 => "001101001",
5408 => "001101000",
5409 => "001100101",
5410 => "001100100",
5411 => "001100110",
5412 => "001100011",
5413 => "001100111",
5414 => "001101101",
5415 => "001101011",
5416 => "001101011",
5417 => "001101010",
5418 => "011100001",
5419 => "010111000",
5420 => "001110001",
5421 => "001100111",
5422 => "001100101",
5423 => "001100101",
5424 => "001100010",
5425 => "001100100",
5426 => "001100011",
5427 => "001100010",
5428 => "001100011",
5429 => "001100011",
5430 => "001100101",
5431 => "001100110",
5432 => "001100110",
5433 => "001100100",
5434 => "001100001",
5435 => "001100011",
5436 => "001011111",
5437 => "001011111",
5438 => "001100011",
5439 => "001100001",
5440 => "001100000",
5441 => "001100010",
5442 => "001011110",
5443 => "001100001",
5444 => "001100001",
5445 => "001100000",
5446 => "001011110",
5447 => "001100000",
5448 => "001100011",
5449 => "001011111",
5450 => "001100000",
5451 => "001100000",
5452 => "001011101",
5453 => "001100000",
5454 => "001100001",
5455 => "001011010",
5456 => "001011100",
5457 => "001011110",
5458 => "001010010",
5459 => "000111101",
5460 => "001000000",
5461 => "000111111",
5462 => "001111100",
5463 => "010111001",
5464 => "011010111",
5465 => "011101100",
5466 => "011010110",
5467 => "011101100",
5468 => "011010110",
5469 => "011011100",
5470 => "010001011",
5471 => "001101000",
5472 => "001100100",
5473 => "001100101",
5474 => "001100101",
5475 => "001100000",
5476 => "001100000",
5477 => "001100001",
5478 => "001100011",
5479 => "001101000",
5480 => "001100100",
5481 => "001100101",
5482 => "001100011",
5483 => "001100100",
5484 => "001100001",
5485 => "001011110",
5486 => "001011101",
5487 => "001100011",
5488 => "001011011",
5489 => "001011011",
5490 => "001011111",
5491 => "001011101",
5492 => "001011100",
5493 => "001100000",
5494 => "001100010",
5495 => "001100001",
5496 => "001100011",
5497 => "001011111",
5498 => "001011110",
5499 => "001011011",
5500 => "001011111",
5501 => "001100001",
5502 => "001011101",
5503 => "001100010",
5504 => "001100000",
5505 => "001100100",
5506 => "001100101",
5507 => "001100100",
5508 => "001100001",
5509 => "001100011",
5510 => "001100101",
5511 => "001100011",
5512 => "001100010",
5513 => "001100011",
5514 => "001100000",
5515 => "001011101",
5516 => "001011110",
5517 => "001011110",
5518 => "001100010",
5519 => "001100011",
5520 => "001100010",
5521 => "001100100",
5522 => "001100011",
5523 => "001100100",
5524 => "001101001",
5525 => "001101010",
5526 => "001100000",
5527 => "001100110",
5528 => "001011110",
5529 => "001100000",
5530 => "001100110",
5531 => "001011111",
5532 => "001100101",
5533 => "001011111",
5534 => "001101001",
5535 => "001100100",
5536 => "001100101",
5537 => "001101000",
5538 => "001101010",
5539 => "001100110",
5540 => "001100101",
5541 => "001100111",
5542 => "001101000",
5543 => "001100111",
5544 => "001100101",
5545 => "010101000",
5546 => "011010000",
5547 => "010000001",
5548 => "001100100",
5549 => "001100101",
5550 => "001100100",
5551 => "001100001",
5552 => "001100101",
5553 => "001100001",
5554 => "001100010",
5555 => "001100010",
5556 => "001100101",
5557 => "001100011",
5558 => "001100010",
5559 => "001100111",
5560 => "001100010",
5561 => "001100001",
5562 => "001100011",
5563 => "001100000",
5564 => "001100000",
5565 => "001100100",
5566 => "001100001",
5567 => "001100011",
5568 => "001100001",
5569 => "001100000",
5570 => "001100000",
5571 => "001100010",
5572 => "001011110",
5573 => "001011111",
5574 => "001011110",
5575 => "001100100",
5576 => "001011110",
5577 => "001100001",
5578 => "001100010",
5579 => "001011110",
5580 => "001100000",
5581 => "001011110",
5582 => "001011100",
5583 => "001011011",
5584 => "001011110",
5585 => "001011010",
5586 => "001010111",
5587 => "001001010",
5588 => "001000110",
5589 => "001000100",
5590 => "010001101",
5591 => "010111000",
5592 => "011100001",
5593 => "011101011",
5594 => "011100101",
5595 => "011101011",
5596 => "011100110",
5597 => "011011110",
5598 => "010001101",
5599 => "001100100",
5600 => "001100110",
5601 => "001101001",
5602 => "001100110",
5603 => "001101010",
5604 => "001101010",
5605 => "001100001",
5606 => "001100101",
5607 => "001011101",
5608 => "001011110",
5609 => "001100001",
5610 => "001100001",
5611 => "001100011",
5612 => "001100011",
5613 => "001100011",
5614 => "001011110",
5615 => "001100101",
5616 => "001100001",
5617 => "001100010",
5618 => "001100010",
5619 => "001100100",
5620 => "001100000",
5621 => "001011101",
5622 => "001011101",
5623 => "001100000",
5624 => "001100001",
5625 => "001011011",
5626 => "001011010",
5627 => "001011110",
5628 => "001100000",
5629 => "001011110",
5630 => "001100001",
5631 => "001100001",
5632 => "001100010",
5633 => "001100000",
5634 => "001100000",
5635 => "001100001",
5636 => "001100101",
5637 => "001100101",
5638 => "001100011",
5639 => "001011110",
5640 => "001100010",
5641 => "001100010",
5642 => "001101000",
5643 => "001100101",
5644 => "001100101",
5645 => "001100111",
5646 => "001101000",
5647 => "001101000",
5648 => "001100000",
5649 => "001100111",
5650 => "001101010",
5651 => "001100011",
5652 => "001100101",
5653 => "001101100",
5654 => "001101001",
5655 => "001101010",
5656 => "001100101",
5657 => "001101001",
5658 => "001100111",
5659 => "001100011",
5660 => "001100100",
5661 => "001100100",
5662 => "001011111",
5663 => "001011010",
5664 => "001011110",
5665 => "001011011",
5666 => "001100001",
5667 => "001011111",
5668 => "001100100",
5669 => "001100010",
5670 => "001101000",
5671 => "001101100",
5672 => "010001001",
5673 => "011001111",
5674 => "010100111",
5675 => "001100111",
5676 => "001100100",
5677 => "001100110",
5678 => "001100100",
5679 => "001100010",
5680 => "001100000",
5681 => "001100011",
5682 => "001100011",
5683 => "001100001",
5684 => "001100011",
5685 => "001100100",
5686 => "001100100",
5687 => "001100110",
5688 => "001100010",
5689 => "001100011",
5690 => "001100000",
5691 => "001100010",
5692 => "001100010",
5693 => "001100010",
5694 => "001011110",
5695 => "001100100",
5696 => "001100010",
5697 => "001011111",
5698 => "001100100",
5699 => "001100000",
5700 => "001100001",
5701 => "001100010",
5702 => "001100000",
5703 => "001011110",
5704 => "001100001",
5705 => "001011101",
5706 => "001011111",
5707 => "001100011",
5708 => "001100000",
5709 => "001011011",
5710 => "001011111",
5711 => "001100010",
5712 => "001011011",
5713 => "001011101",
5714 => "001011100",
5715 => "001011001",
5716 => "001001010",
5717 => "001000110",
5718 => "010100110",
5719 => "011000001",
5720 => "011011100",
5721 => "011100111",
5722 => "011110000",
5723 => "011110001",
5724 => "011100010",
5725 => "011101010",
5726 => "010000111",
5727 => "001100100",
5728 => "001100010",
5729 => "001101100",
5730 => "001100011",
5731 => "001100101",
5732 => "001011101",
5733 => "001100100",
5734 => "001101001",
5735 => "001100110",
5736 => "001100110",
5737 => "001100011",
5738 => "001100100",
5739 => "001100010",
5740 => "001100110",
5741 => "001100101",
5742 => "001100010",
5743 => "001100011",
5744 => "001100100",
5745 => "001100011",
5746 => "001100011",
5747 => "001100000",
5748 => "001011100",
5749 => "001011111",
5750 => "001011111",
5751 => "001011111",
5752 => "001011001",
5753 => "001011010",
5754 => "001100000",
5755 => "001100001",
5756 => "001100001",
5757 => "001100000",
5758 => "001100000",
5759 => "001100000",
5760 => "001011101",
5761 => "001011101",
5762 => "001010111",
5763 => "001010110",
5764 => "001010110",
5765 => "001011011",
5766 => "001100010",
5767 => "001100001",
5768 => "001100110",
5769 => "001100110",
5770 => "001100110",
5771 => "001100101",
5772 => "001101001",
5773 => "001100110",
5774 => "001100111",
5775 => "001101000",
5776 => "001100111",
5777 => "001100111",
5778 => "001101010",
5779 => "001101000",
5780 => "001101000",
5781 => "001100110",
5782 => "001100011",
5783 => "001100100",
5784 => "001101001",
5785 => "001100111",
5786 => "001100101",
5787 => "001100101",
5788 => "001100111",
5789 => "001100100",
5790 => "001100011",
5791 => "001100011",
5792 => "001100100",
5793 => "001100100",
5794 => "001100101",
5795 => "001100100",
5796 => "001100110",
5797 => "001101001",
5798 => "001100101",
5799 => "001111010",
5800 => "011011010",
5801 => "010101100",
5802 => "001100111",
5803 => "001100100",
5804 => "001100100",
5805 => "001100101",
5806 => "001100100",
5807 => "001100100",
5808 => "001100010",
5809 => "001100100",
5810 => "001100011",
5811 => "001100011",
5812 => "001100011",
5813 => "001100000",
5814 => "001100010",
5815 => "001100010",
5816 => "001100100",
5817 => "001100001",
5818 => "001100000",
5819 => "001100100",
5820 => "001100011",
5821 => "001011111",
5822 => "001100010",
5823 => "001100001",
5824 => "001100001",
5825 => "001100100",
5826 => "001100010",
5827 => "001100001",
5828 => "001100010",
5829 => "001100001",
5830 => "001100010",
5831 => "001100011",
5832 => "001100000",
5833 => "001011110",
5834 => "001100010",
5835 => "001011111",
5836 => "001011110",
5837 => "001100000",
5838 => "001011111",
5839 => "001011110",
5840 => "001011111",
5841 => "001011111",
5842 => "001011110",
5843 => "001011011",
5844 => "001011100",
5845 => "001010001",
5846 => "010101001",
5847 => "011000011",
5848 => "011011010",
5849 => "011110001",
5850 => "011101001",
5851 => "011011110",
5852 => "011100010",
5853 => "011110011",
5854 => "011011110",
5855 => "001101101",
5856 => "001101101",
5857 => "001101001",
5858 => "001100011",
5859 => "001100111",
5860 => "001100111",
5861 => "001100110",
5862 => "001100111",
5863 => "001100110",
5864 => "001100101",
5865 => "001101000",
5866 => "001101000",
5867 => "001100101",
5868 => "001011110",
5869 => "001100000",
5870 => "001011111",
5871 => "001100001",
5872 => "001011110",
5873 => "001011111",
5874 => "001100000",
5875 => "001011101",
5876 => "001011100",
5877 => "001011110",
5878 => "001011110",
5879 => "001100001",
5880 => "001100011",
5881 => "001011110",
5882 => "001011100",
5883 => "001100011",
5884 => "001100000",
5885 => "001100011",
5886 => "001100011",
5887 => "001011111",
5888 => "001011111",
5889 => "001011110",
5890 => "001011100",
5891 => "001100000",
5892 => "001011100",
5893 => "001100010",
5894 => "001011111",
5895 => "001011111",
5896 => "001011111",
5897 => "001011111",
5898 => "001100001",
5899 => "001100011",
5900 => "001100011",
5901 => "001100100",
5902 => "001100100",
5903 => "001100000",
5904 => "001100100",
5905 => "001100111",
5906 => "001101010",
5907 => "001100111",
5908 => "001100100",
5909 => "001101000",
5910 => "001101000",
5911 => "001101011",
5912 => "001101010",
5913 => "001101000",
5914 => "001100101",
5915 => "001100101",
5916 => "001100010",
5917 => "001100011",
5918 => "001100011",
5919 => "001100110",
5920 => "001101000",
5921 => "001101001",
5922 => "001100110",
5923 => "001100011",
5924 => "001100100",
5925 => "001100110",
5926 => "001101111",
5927 => "011000110",
5928 => "010111100",
5929 => "001101000",
5930 => "001100110",
5931 => "001100010",
5932 => "001100001",
5933 => "001100010",
5934 => "001100011",
5935 => "001011111",
5936 => "001100011",
5937 => "001100001",
5938 => "001100001",
5939 => "001100000",
5940 => "001100001",
5941 => "001100011",
5942 => "001100011",
5943 => "001100100",
5944 => "001100010",
5945 => "001100000",
5946 => "001100001",
5947 => "001100000",
5948 => "001100001",
5949 => "001100010",
5950 => "001100001",
5951 => "001100011",
5952 => "001100101",
5953 => "001100011",
5954 => "001100000",
5955 => "001100010",
5956 => "001100011",
5957 => "001100001",
5958 => "001100000",
5959 => "001011111",
5960 => "001011110",
5961 => "001101000",
5962 => "001011110",
5963 => "001011111",
5964 => "001011111",
5965 => "001011110",
5966 => "001100000",
5967 => "001011111",
5968 => "001100010",
5969 => "001100010",
5970 => "001100011",
5971 => "001100001",
5972 => "001100001",
5973 => "001101010",
5974 => "010111001",
5975 => "011100101",
5976 => "011110000",
5977 => "011101000",
5978 => "011101011",
5979 => "011101110",
5980 => "011101001",
5981 => "011110011",
5982 => "011101000",
5983 => "011000000",
5984 => "001101011",
5985 => "001100110",
5986 => "001100101",
5987 => "001100100",
5988 => "001100100",
5989 => "001100010",
5990 => "001100110",
5991 => "001100011",
5992 => "001100011",
5993 => "001100101",
5994 => "001100001",
5995 => "001100000",
5996 => "001100011",
5997 => "001100001",
5998 => "001100010",
5999 => "001100001",
6000 => "001011111",
6001 => "001011100",
6002 => "001100001",
6003 => "001011110",
6004 => "001011101",
6005 => "001011010",
6006 => "001011000",
6007 => "001010111",
6008 => "001011100",
6009 => "001011110",
6010 => "001011110",
6011 => "001011100",
6012 => "001011101",
6013 => "001011111",
6014 => "001011110",
6015 => "001011011",
6016 => "001011111",
6017 => "001011110",
6018 => "001100010",
6019 => "001100010",
6020 => "001100000",
6021 => "001100010",
6022 => "001100010",
6023 => "001100001",
6024 => "001100010",
6025 => "001100001",
6026 => "001011110",
6027 => "001011101",
6028 => "001100000",
6029 => "001100110",
6030 => "001100101",
6031 => "001011111",
6032 => "001011111",
6033 => "001101100",
6034 => "001100011",
6035 => "001100011",
6036 => "001100001",
6037 => "001100011",
6038 => "001100100",
6039 => "001100101",
6040 => "001100101",
6041 => "001100111",
6042 => "001100111",
6043 => "001101111",
6044 => "001110011",
6045 => "001111000",
6046 => "001111100",
6047 => "010000010",
6048 => "001110101",
6049 => "001111001",
6050 => "001110100",
6051 => "001101110",
6052 => "001110000",
6053 => "001101111",
6054 => "010011011",
6055 => "011000100",
6056 => "001101011",
6057 => "001100010",
6058 => "001100010",
6059 => "001100011",
6060 => "001100011",
6061 => "001100010",
6062 => "001100001",
6063 => "001100011",
6064 => "001100011",
6065 => "001100011",
6066 => "001100100",
6067 => "001100001",
6068 => "001100011",
6069 => "001100011",
6070 => "001100010",
6071 => "001100010",
6072 => "001100010",
6073 => "001100011",
6074 => "001100000",
6075 => "001100001",
6076 => "001100010",
6077 => "001100010",
6078 => "001100000",
6079 => "001100010",
6080 => "001100000",
6081 => "001100011",
6082 => "001100101",
6083 => "001100001",
6084 => "001100000",
6085 => "001100001",
6086 => "001100001",
6087 => "001100000",
6088 => "001100011",
6089 => "001011111",
6090 => "001100000",
6091 => "001100001",
6092 => "001011111",
6093 => "001100000",
6094 => "001100000",
6095 => "001011111",
6096 => "001100010",
6097 => "001100001",
6098 => "001011110",
6099 => "001100000",
6100 => "001100101",
6101 => "010010011",
6102 => "011011101",
6103 => "011110011",
6104 => "011101101",
6105 => "011101001",
6106 => "011100001",
6107 => "011100101",
6108 => "011100101",
6109 => "011101111",
6110 => "011011001",
6111 => "011011101",
6112 => "010011100",
6113 => "001101010",
6114 => "001101100",
6115 => "001100111",
6116 => "001100101",
6117 => "001100011",
6118 => "001100101",
6119 => "001100000",
6120 => "001100001",
6121 => "001100000",
6122 => "001011111",
6123 => "001100000",
6124 => "001100001",
6125 => "001011101",
6126 => "001011100",
6127 => "001011011",
6128 => "001011111",
6129 => "001011101",
6130 => "001011110",
6131 => "001011101",
6132 => "001011011",
6133 => "001011011",
6134 => "001011001",
6135 => "001011000",
6136 => "001011011",
6137 => "001011001",
6138 => "001011101",
6139 => "001011101",
6140 => "001011011",
6141 => "001011101",
6142 => "001011100",
6143 => "001011100",
6144 => "001100000",
6145 => "001100001",
6146 => "001011101",
6147 => "001011000",
6148 => "001100000",
6149 => "001101010",
6150 => "001101101",
6151 => "001110000",
6152 => "001101111",
6153 => "001110000",
6154 => "001101110",
6155 => "001111101",
6156 => "010000010",
6157 => "001111000",
6158 => "001111001",
6159 => "001111010",
6160 => "001101011",
6161 => "001101101",
6162 => "001101100",
6163 => "010000001",
6164 => "001110110",
6165 => "010000010",
6166 => "001111001",
6167 => "001111011",
6168 => "001110101",
6169 => "001110001",
6170 => "001111101",
6171 => "001101111",
6172 => "001101111",
6173 => "001101110",
6174 => "001101010",
6175 => "001101010",
6176 => "001111011",
6177 => "001110010",
6178 => "001110001",
6179 => "001110001",
6180 => "001111001",
6181 => "001111011",
6182 => "010010111",
6183 => "001101000",
6184 => "001100011",
6185 => "001100010",
6186 => "001100111",
6187 => "001100110",
6188 => "001100011",
6189 => "001100001",
6190 => "001100100",
6191 => "001100101",
6192 => "001100011",
6193 => "001100011",
6194 => "001100011",
6195 => "001100000",
6196 => "001100011",
6197 => "001100001",
6198 => "001100011",
6199 => "001100011",
6200 => "001100011",
6201 => "001100011",
6202 => "001011111",
6203 => "001100001",
6204 => "001100000",
6205 => "001100001",
6206 => "001100011",
6207 => "001100010",
6208 => "001100000",
6209 => "001100011",
6210 => "001100001",
6211 => "001100100",
6212 => "001100011",
6213 => "001100010",
6214 => "001011111",
6215 => "001100000",
6216 => "001100000",
6217 => "001100010",
6218 => "001100010",
6219 => "001100000",
6220 => "001100000",
6221 => "001100011",
6222 => "001100001",
6223 => "001100010",
6224 => "001100010",
6225 => "001011111",
6226 => "001100010",
6227 => "001100110",
6228 => "001110110",
6229 => "011010000",
6230 => "011101111",
6231 => "011110010",
6232 => "011110000",
6233 => "011101100",
6234 => "011101011",
6235 => "011101111",
6236 => "011100001",
6237 => "011100111",
6238 => "011100010",
6239 => "011100011",
6240 => "011101000",
6241 => "010001101",
6242 => "001101000",
6243 => "001100101",
6244 => "001100011",
6245 => "001100101",
6246 => "001100001",
6247 => "001011101",
6248 => "001100011",
6249 => "001011101",
6250 => "001011110",
6251 => "001011111",
6252 => "001011110",
6253 => "001100011",
6254 => "001101010",
6255 => "001100000",
6256 => "001100000",
6257 => "001100010",
6258 => "001100001",
6259 => "001100001",
6260 => "001100010",
6261 => "001100000",
6262 => "001100001",
6263 => "001100100",
6264 => "001100000",
6265 => "001100001",
6266 => "001011111",
6267 => "001011111",
6268 => "001011111",
6269 => "001011011",
6270 => "001011011",
6271 => "001011101",
6272 => "001111011",
6273 => "001111010",
6274 => "000111100",
6275 => "001001111",
6276 => "001011100",
6277 => "001110001",
6278 => "001101110",
6279 => "001101010",
6280 => "001100110",
6281 => "001100101",
6282 => "001110100",
6283 => "010010111",
6284 => "010010110",
6285 => "001101000",
6286 => "001100001",
6287 => "001101101",
6288 => "001101010",
6289 => "001101110",
6290 => "001110000",
6291 => "001111101",
6292 => "001101100",
6293 => "010001110",
6294 => "010001100",
6295 => "001110100",
6296 => "001110111",
6297 => "001101110",
6298 => "001111001",
6299 => "001110000",
6300 => "001111001",
6301 => "001100100",
6302 => "001011111",
6303 => "001100100",
6304 => "001110000",
6305 => "001011011",
6306 => "001100111",
6307 => "001110111",
6308 => "001001111",
6309 => "001001011",
6310 => "010000000",
6311 => "010000100",
6312 => "001110011",
6313 => "001100011",
6314 => "001011001",
6315 => "001010111",
6316 => "001100101",
6317 => "001100011",
6318 => "001100110",
6319 => "001100011",
6320 => "001100001",
6321 => "001100011",
6322 => "001100000",
6323 => "001100100",
6324 => "001100100",
6325 => "001100011",
6326 => "001100001",
6327 => "001100010",
6328 => "001100010",
6329 => "001100010",
6330 => "001100001",
6331 => "001100100",
6332 => "001100011",
6333 => "001100011",
6334 => "001100010",
6335 => "001100100",
6336 => "001100100",
6337 => "001100010",
6338 => "001100010",
6339 => "001100011",
6340 => "001100000",
6341 => "001100000",
6342 => "001100000",
6343 => "001011110",
6344 => "001100010",
6345 => "001100001",
6346 => "001011111",
6347 => "001011111",
6348 => "001100010",
6349 => "001100011",
6350 => "001100010",
6351 => "001100001",
6352 => "001100010",
6353 => "001100010",
6354 => "001101000",
6355 => "001101100",
6356 => "011011011",
6357 => "011101101",
6358 => "011110101",
6359 => "011110001",
6360 => "011110001",
6361 => "011101101",
6362 => "011101011",
6363 => "011101101",
6364 => "011101110",
6365 => "011110100",
6366 => "011110101",
6367 => "011110101",
6368 => "011100010",
6369 => "011100100",
6370 => "010000010",
6371 => "001101001",
6372 => "001100101",
6373 => "001100110",
6374 => "001100110",
6375 => "001100111",
6376 => "001100111",
6377 => "001100101",
6378 => "001100100",
6379 => "001100010",
6380 => "001100110",
6381 => "001100101",
6382 => "001100011",
6383 => "001100011",
6384 => "001100110",
6385 => "001100100",
6386 => "001100010",
6387 => "001011111",
6388 => "001100000",
6389 => "001100001",
6390 => "001100000",
6391 => "001100011",
6392 => "001100111",
6393 => "001100011",
6394 => "001011100",
6395 => "001011000",
6396 => "001011110",
6397 => "001011101",
6398 => "001011101",
6399 => "001011001",
6400 => "001100101",
6401 => "001101000",
6402 => "000111011",
6403 => "001001000",
6404 => "001100001",
6405 => "001101101",
6406 => "001101011",
6407 => "001101010",
6408 => "001101110",
6409 => "001101010",
6410 => "001111010",
6411 => "010010001",
6412 => "010010000",
6413 => "001110001",
6414 => "001110000",
6415 => "001010101",
6416 => "001101001",
6417 => "001101100",
6418 => "001101011",
6419 => "001101010",
6420 => "001100010",
6421 => "010010000",
6422 => "010001000",
6423 => "001100111",
6424 => "001010100",
6425 => "001000111",
6426 => "001011010",
6427 => "001000111",
6428 => "001110000",
6429 => "001100010",
6430 => "001001110",
6431 => "001010000",
6432 => "001100000",
6433 => "001010110",
6434 => "001101011",
6435 => "001110000",
6436 => "001001101",
6437 => "001001010",
6438 => "010000011",
6439 => "010110000",
6440 => "010101111",
6441 => "010100111",
6442 => "010011111",
6443 => "010001001",
6444 => "001101101",
6445 => "001011111",
6446 => "001011100",
6447 => "001011100",
6448 => "001100001",
6449 => "001100010",
6450 => "001100011",
6451 => "001100001",
6452 => "001011111",
6453 => "001100100",
6454 => "001100001",
6455 => "001100001",
6456 => "001100001",
6457 => "001100001",
6458 => "001100001",
6459 => "001100000",
6460 => "001100010",
6461 => "001100011",
6462 => "001100011",
6463 => "001100100",
6464 => "001100001",
6465 => "001100100",
6466 => "001100011",
6467 => "001100000",
6468 => "001100101",
6469 => "001100001",
6470 => "001011111",
6471 => "001100011",
6472 => "001100010",
6473 => "001100000",
6474 => "001100000",
6475 => "001011111",
6476 => "001100010",
6477 => "001100100",
6478 => "001100001",
6479 => "001100000",
6480 => "001100001",
6481 => "001100111",
6482 => "001101011",
6483 => "011001111",
6484 => "011101000",
6485 => "011101000",
6486 => "011110101",
6487 => "011110001",
6488 => "011110100",
6489 => "011110001",
6490 => "011110000",
6491 => "011101111",
6492 => "011101100",
6493 => "011100100",
6494 => "011101001",
6495 => "011100101",
6496 => "011100110",
6497 => "011100011",
6498 => "011001110",
6499 => "001111001",
6500 => "001101110",
6501 => "001101001",
6502 => "001101000",
6503 => "001101101",
6504 => "001101101",
6505 => "001101100",
6506 => "001101010",
6507 => "001100101",
6508 => "001101000",
6509 => "001100110",
6510 => "001100110",
6511 => "001100010",
6512 => "001100100",
6513 => "001100100",
6514 => "001100100",
6515 => "001100000",
6516 => "001100010",
6517 => "001100100",
6518 => "001100001",
6519 => "001100010",
6520 => "001100011",
6521 => "001100010",
6522 => "001100011",
6523 => "001100011",
6524 => "001100000",
6525 => "001011111",
6526 => "001011111",
6527 => "001100001",
6528 => "001001010",
6529 => "000111000",
6530 => "001000000",
6531 => "001000001",
6532 => "001000110",
6533 => "001000010",
6534 => "001000101",
6535 => "000111111",
6536 => "001000110",
6537 => "000111110",
6538 => "001010101",
6539 => "010010010",
6540 => "010001000",
6541 => "001001001",
6542 => "000111000",
6543 => "000101110",
6544 => "001100000",
6545 => "001101001",
6546 => "001100001",
6547 => "001000001",
6548 => "000110100",
6549 => "010010111",
6550 => "010010000",
6551 => "010000101",
6552 => "001010110",
6553 => "001011100",
6554 => "001010011",
6555 => "001001110",
6556 => "001110011",
6557 => "001101000",
6558 => "001101011",
6559 => "001010110",
6560 => "001010110",
6561 => "001000111",
6562 => "001100110",
6563 => "001001100",
6564 => "001001000",
6565 => "000111110",
6566 => "010001001",
6567 => "010111111",
6568 => "011001001",
6569 => "011000010",
6570 => "011000000",
6571 => "010101100",
6572 => "010100110",
6573 => "010100011",
6574 => "010011011",
6575 => "010000011",
6576 => "001011110",
6577 => "001100010",
6578 => "001100010",
6579 => "001100100",
6580 => "001100100",
6581 => "001100011",
6582 => "001100011",
6583 => "001011111",
6584 => "001100001",
6585 => "001100010",
6586 => "001100001",
6587 => "001100100",
6588 => "001100010",
6589 => "001100001",
6590 => "001100000",
6591 => "001100010",
6592 => "001100100",
6593 => "001100001",
6594 => "001100010",
6595 => "001100011",
6596 => "001100001",
6597 => "001100001",
6598 => "001100010",
6599 => "001011111",
6600 => "001100001",
6601 => "001100011",
6602 => "001100010",
6603 => "001100001",
6604 => "001100010",
6605 => "001100001",
6606 => "001100001",
6607 => "001100100",
6608 => "001100011",
6609 => "001100110",
6610 => "010101000",
6611 => "011010101",
6612 => "011110010",
6613 => "011110110",
6614 => "011110101",
6615 => "011110100",
6616 => "011110101",
6617 => "011110100",
6618 => "011110010",
6619 => "011101111",
6620 => "011110001",
6621 => "011101001",
6622 => "011101100",
6623 => "011100101",
6624 => "011100010",
6625 => "011101110",
6626 => "011101110",
6627 => "011010101",
6628 => "001110111",
6629 => "001110001",
6630 => "001110000",
6631 => "001110000",
6632 => "001110000",
6633 => "001101101",
6634 => "001110000",
6635 => "001101101",
6636 => "001101110",
6637 => "001101011",
6638 => "001101000",
6639 => "001101001",
6640 => "001100100",
6641 => "001101010",
6642 => "001101001",
6643 => "001101010",
6644 => "001101000",
6645 => "001100111",
6646 => "001101010",
6647 => "001101011",
6648 => "001101001",
6649 => "001101000",
6650 => "001100110",
6651 => "001100111",
6652 => "001100111",
6653 => "001100100",
6654 => "001100100",
6655 => "001100011",
6656 => "001000111",
6657 => "000110110",
6658 => "001000010",
6659 => "001000010",
6660 => "001011011",
6661 => "001011111",
6662 => "001100010",
6663 => "001011101",
6664 => "001010101",
6665 => "001000001",
6666 => "001010101",
6667 => "010001110",
6668 => "010000011",
6669 => "001011000",
6670 => "001010111",
6671 => "000111100",
6672 => "001100010",
6673 => "001100111",
6674 => "001100011",
6675 => "001010100",
6676 => "000110100",
6677 => "010000101",
6678 => "010010101",
6679 => "010001000",
6680 => "001010110",
6681 => "001010011",
6682 => "001010111",
6683 => "000111101",
6684 => "001101000",
6685 => "001101011",
6686 => "001100111",
6687 => "001011000",
6688 => "001010110",
6689 => "001010001",
6690 => "001000011",
6691 => "001001000",
6692 => "000111111",
6693 => "000111111",
6694 => "010001100",
6695 => "011000010",
6696 => "011000100",
6697 => "011000101",
6698 => "011000110",
6699 => "011000010",
6700 => "010111110",
6701 => "011000001",
6702 => "010001111",
6703 => "001100101",
6704 => "001100011",
6705 => "001100100",
6706 => "001100100",
6707 => "001100011",
6708 => "001100011",
6709 => "001100100",
6710 => "001100001",
6711 => "001100010",
6712 => "001100011",
6713 => "001100101",
6714 => "001100011",
6715 => "001100101",
6716 => "001100011",
6717 => "001100010",
6718 => "001100100",
6719 => "001100010",
6720 => "001100010",
6721 => "001100001",
6722 => "001100100",
6723 => "001100000",
6724 => "001100001",
6725 => "001100110",
6726 => "001011111",
6727 => "001100001",
6728 => "001100100",
6729 => "001100001",
6730 => "001100010",
6731 => "001100011",
6732 => "001100010",
6733 => "001100001",
6734 => "001100001",
6735 => "001100011",
6736 => "001100111",
6737 => "010000100",
6738 => "011010111",
6739 => "011100100",
6740 => "011110100",
6741 => "011110110",
6742 => "011101111",
6743 => "011110010",
6744 => "011110011",
6745 => "011110101",
6746 => "011110101",
6747 => "011101101",
6748 => "011110000",
6749 => "011110100",
6750 => "011110001",
6751 => "011101011",
6752 => "011101010",
6753 => "011101000",
6754 => "011101101",
6755 => "011101100",
6756 => "011010011",
6757 => "001100111",
6758 => "001100110",
6759 => "001100011",
6760 => "001011101",
6761 => "001100011",
6762 => "001100000",
6763 => "001100010",
6764 => "001011110",
6765 => "001100110",
6766 => "001100110",
6767 => "001100010",
6768 => "001100100",
6769 => "001100100",
6770 => "001100011",
6771 => "001100100",
6772 => "001100101",
6773 => "001100011",
6774 => "001100011",
6775 => "001100101",
6776 => "001101000",
6777 => "001101000",
6778 => "001101001",
6779 => "001101010",
6780 => "001101101",
6781 => "001101010",
6782 => "001101001",
6783 => "001101000",
6784 => "001011101",
6785 => "001000001",
6786 => "001000011",
6787 => "001000010",
6788 => "001001111",
6789 => "001011100",
6790 => "001100101",
6791 => "001011010",
6792 => "001011110",
6793 => "001010001",
6794 => "001011111",
6795 => "001110111",
6796 => "001111010",
6797 => "001010101",
6798 => "001011101",
6799 => "001011001",
6800 => "001100110",
6801 => "001101010",
6802 => "001100011",
6803 => "001011100",
6804 => "001010001",
6805 => "001010111",
6806 => "001100100",
6807 => "001011100",
6808 => "001011011",
6809 => "001011000",
6810 => "001011000",
6811 => "001011011",
6812 => "001010110",
6813 => "001010111",
6814 => "001011011",
6815 => "001011011",
6816 => "001011001",
6817 => "000111100",
6818 => "000111100",
6819 => "000110010",
6820 => "000110111",
6821 => "000111010",
6822 => "010010001",
6823 => "011000100",
6824 => "010111111",
6825 => "011000100",
6826 => "011000101",
6827 => "011000010",
6828 => "010111101",
6829 => "011000011",
6830 => "001010110",
6831 => "001010110",
6832 => "001011011",
6833 => "001100110",
6834 => "001100100",
6835 => "001100100",
6836 => "001100101",
6837 => "001100100",
6838 => "001100101",
6839 => "001100011",
6840 => "001100011",
6841 => "001010011",
6842 => "001011100",
6843 => "001100100",
6844 => "001100011",
6845 => "001100011",
6846 => "001100011",
6847 => "001100010",
6848 => "001100010",
6849 => "001100010",
6850 => "001100001",
6851 => "001100001",
6852 => "001100001",
6853 => "001100000",
6854 => "001100010",
6855 => "001100011",
6856 => "001100011",
6857 => "001100100",
6858 => "001100000",
6859 => "001100000",
6860 => "001100010",
6861 => "001100001",
6862 => "001100011",
6863 => "001100110",
6864 => "001111011",
6865 => "011011010",
6866 => "011100011",
6867 => "011110100",
6868 => "011110101",
6869 => "011110101",
6870 => "011110100",
6871 => "011110010",
6872 => "011110110",
6873 => "011110101",
6874 => "011110110",
6875 => "011110000",
6876 => "011110101",
6877 => "011110110",
6878 => "011110010",
6879 => "011100111",
6880 => "011100000",
6881 => "011011101",
6882 => "011101001",
6883 => "011110010",
6884 => "011110000",
6885 => "010110110",
6886 => "001100010",
6887 => "001100001",
6888 => "001100011",
6889 => "001100100",
6890 => "001101011",
6891 => "001100110",
6892 => "001100100",
6893 => "001100100",
6894 => "001100010",
6895 => "001100001",
6896 => "001100011",
6897 => "001100010",
6898 => "001100010",
6899 => "001100011",
6900 => "001100010",
6901 => "001100100",
6902 => "001100100",
6903 => "001100001",
6904 => "001100101",
6905 => "001100101",
6906 => "001100011",
6907 => "001100111",
6908 => "001100111",
6909 => "001100111",
6910 => "001101001",
6911 => "001100101",
6912 => "001100001",
6913 => "001010110",
6914 => "001011001",
6915 => "001011101",
6916 => "001011010",
6917 => "001011110",
6918 => "001011101",
6919 => "001011101",
6920 => "001100000",
6921 => "001100001",
6922 => "001100011",
6923 => "001100001",
6924 => "001011111",
6925 => "001011001",
6926 => "001010100",
6927 => "001010011",
6928 => "001100000",
6929 => "001100000",
6930 => "001011110",
6931 => "001011111",
6932 => "001100001",
6933 => "001011100",
6934 => "001011101",
6935 => "001011100",
6936 => "001100010",
6937 => "001011011",
6938 => "001011110",
6939 => "001011110",
6940 => "001011101",
6941 => "001011001",
6942 => "001011010",
6943 => "001011010",
6944 => "001001011",
6945 => "000111111",
6946 => "001001001",
6947 => "000110000",
6948 => "000110101",
6949 => "001000000",
6950 => "010010011",
6951 => "011000000",
6952 => "011000010",
6953 => "011001000",
6954 => "011000100",
6955 => "011000111",
6956 => "010111101",
6957 => "010101100",
6958 => "001101111",
6959 => "010101001",
6960 => "010100001",
6961 => "010010100",
6962 => "001110011",
6963 => "001010001",
6964 => "001011010",
6965 => "001100111",
6966 => "001100100",
6967 => "001100110",
6968 => "010101010",
6969 => "010110100",
6970 => "010100111",
6971 => "010011101",
6972 => "001111110",
6973 => "001011100",
6974 => "001011000",
6975 => "001100011",
6976 => "001100110",
6977 => "001100010",
6978 => "001100000",
6979 => "001100010",
6980 => "001100001",
6981 => "001100100",
6982 => "001100010",
6983 => "001100001",
6984 => "001100011",
6985 => "001100011",
6986 => "001100010",
6987 => "001100010",
6988 => "001100001",
6989 => "001100011",
6990 => "001101000",
6991 => "001101110",
6992 => "011010000",
6993 => "011010011",
6994 => "011110100",
6995 => "011110101",
6996 => "011110011",
6997 => "011110011",
6998 => "011110011",
6999 => "011110011",
7000 => "011110011",
7001 => "011110110",
7002 => "011110011",
7003 => "011101111",
7004 => "011110001",
7005 => "011110010",
7006 => "011110101",
7007 => "011110011",
7008 => "011110010",
7009 => "011101111",
7010 => "011101100",
7011 => "011101001",
7012 => "011110011",
7013 => "011101010",
7014 => "001010001",
7015 => "001001111",
7016 => "001001110",
7017 => "001001101",
7018 => "001010010",
7019 => "001001110",
7020 => "001011011",
7021 => "001011000",
7022 => "001100100",
7023 => "001101001",
7024 => "001101001",
7025 => "001100110",
7026 => "001100011",
7027 => "001100010",
7028 => "001100000",
7029 => "001100010",
7030 => "001100000",
7031 => "001011111",
7032 => "001011111",
7033 => "001011100",
7034 => "001011110",
7035 => "001011100",
7036 => "001011101",
7037 => "001011111",
7038 => "001100011",
7039 => "001100001",
7040 => "001110001",
7041 => "001101110",
7042 => "001100101",
7043 => "001100100",
7044 => "001100110",
7045 => "001100011",
7046 => "001100100",
7047 => "001100101",
7048 => "001011111",
7049 => "001011101",
7050 => "001011101",
7051 => "001011110",
7052 => "001011111",
7053 => "001100000",
7054 => "001011110",
7055 => "001011111",
7056 => "001100000",
7057 => "001011111",
7058 => "001011110",
7059 => "001100001",
7060 => "001100011",
7061 => "001100000",
7062 => "001100010",
7063 => "001100011",
7064 => "001100100",
7065 => "001100010",
7066 => "001101100",
7067 => "001101010",
7068 => "001100011",
7069 => "001100010",
7070 => "001100001",
7071 => "001011010",
7072 => "001010001",
7073 => "001001001",
7074 => "011011111",
7075 => "010000011",
7076 => "000101101",
7077 => "000101110",
7078 => "010010111",
7079 => "010111111",
7080 => "010111111",
7081 => "011000010",
7082 => "011000101",
7083 => "010110110",
7084 => "010101101",
7085 => "010011110",
7086 => "001111101",
7087 => "011000010",
7088 => "011000100",
7089 => "010111001",
7090 => "010101110",
7091 => "010100101",
7092 => "010011100",
7093 => "010001101",
7094 => "001101011",
7095 => "011000001",
7096 => "011101001",
7097 => "011110001",
7098 => "010111101",
7099 => "010110100",
7100 => "010101000",
7101 => "010100000",
7102 => "010011010",
7103 => "010001101",
7104 => "001111010",
7105 => "001011011",
7106 => "001010101",
7107 => "001100011",
7108 => "001100011",
7109 => "001100010",
7110 => "001100001",
7111 => "001100100",
7112 => "001100001",
7113 => "001100000",
7114 => "001100100",
7115 => "001100001",
7116 => "001100000",
7117 => "001100110",
7118 => "001100011",
7119 => "011000111",
7120 => "011001110",
7121 => "011110000",
7122 => "011110011",
7123 => "011110000",
7124 => "011110011",
7125 => "011110100",
7126 => "011110110",
7127 => "011110100",
7128 => "011110110",
7129 => "011110110",
7130 => "011110000",
7131 => "011110010",
7132 => "011101111",
7133 => "011110110",
7134 => "011101110",
7135 => "011110010",
7136 => "011101110",
7137 => "011101110",
7138 => "011101100",
7139 => "011100111",
7140 => "011101001",
7141 => "011010110",
7142 => "001010001",
7143 => "001010000",
7144 => "001010001",
7145 => "001001111",
7146 => "001001101",
7147 => "001001011",
7148 => "001001101",
7149 => "001001100",
7150 => "001010001",
7151 => "001011100",
7152 => "001011100",
7153 => "001011111",
7154 => "010000100",
7155 => "001110010",
7156 => "001100100",
7157 => "001100001",
7158 => "001100010",
7159 => "001100010",
7160 => "001011111",
7161 => "001100000",
7162 => "001011111",
7163 => "001100001",
7164 => "001100000",
7165 => "001011111",
7166 => "001100001",
7167 => "001100001",
7168 => "001101100",
7169 => "001011010",
7170 => "001011110",
7171 => "001100011",
7172 => "001100100",
7173 => "001100001",
7174 => "001011011",
7175 => "001100111",
7176 => "001101001",
7177 => "001101101",
7178 => "001101111",
7179 => "001101001",
7180 => "001101011",
7181 => "001101111",
7182 => "001100010",
7183 => "001101011",
7184 => "001100100",
7185 => "001100100",
7186 => "001100100",
7187 => "001100100",
7188 => "001100100",
7189 => "001100101",
7190 => "001100010",
7191 => "001100100",
7192 => "001100110",
7193 => "001100110",
7194 => "001100000",
7195 => "001100111",
7196 => "001100100",
7197 => "001011110",
7198 => "001100111",
7199 => "001100011",
7200 => "001100001",
7201 => "010110100",
7202 => "011101010",
7203 => "011110011",
7204 => "001000000",
7205 => "000110100",
7206 => "010010111",
7207 => "010110110",
7208 => "010110110",
7209 => "010111011",
7210 => "011000011",
7211 => "010101011",
7212 => "010100111",
7213 => "010011100",
7214 => "001111110",
7215 => "011000101",
7216 => "011000101",
7217 => "011000001",
7218 => "011000110",
7219 => "011000001",
7220 => "010111110",
7221 => "010110010",
7222 => "010111110",
7223 => "011100111",
7224 => "011110000",
7225 => "011110101",
7226 => "011010000",
7227 => "011000100",
7228 => "011000000",
7229 => "010110011",
7230 => "010101000",
7231 => "010100000",
7232 => "010100000",
7233 => "010011100",
7234 => "010010100",
7235 => "010000110",
7236 => "001110110",
7237 => "001011110",
7238 => "001010100",
7239 => "001011111",
7240 => "001100000",
7241 => "001100100",
7242 => "001100001",
7243 => "001100100",
7244 => "001100111",
7245 => "001100011",
7246 => "010110011",
7247 => "011010010",
7248 => "011011011",
7249 => "011110011",
7250 => "011110011",
7251 => "011110010",
7252 => "011110101",
7253 => "011101010",
7254 => "011110010",
7255 => "011110101",
7256 => "011110101",
7257 => "011110101",
7258 => "011101110",
7259 => "011110011",
7260 => "011110011",
7261 => "011110101",
7262 => "011110100",
7263 => "011101111",
7264 => "011101100",
7265 => "011110010",
7266 => "011110001",
7267 => "011110011",
7268 => "010111000",
7269 => "011010100",
7270 => "001010101",
7271 => "001010010",
7272 => "001001111",
7273 => "001001111",
7274 => "001001101",
7275 => "001001110",
7276 => "001001111",
7277 => "001001010",
7278 => "001011100",
7279 => "011010011",
7280 => "011011110",
7281 => "010100011",
7282 => "011110011",
7283 => "011010011",
7284 => "001011110",
7285 => "001011111",
7286 => "001100000",
7287 => "001100001",
7288 => "001011111",
7289 => "001100100",
7290 => "001101011",
7291 => "001101010",
7292 => "001101010",
7293 => "001011100",
7294 => "001011011",
7295 => "001011100",
7296 => "001011011",
7297 => "001100100",
7298 => "001100111",
7299 => "001100111",
7300 => "001100010",
7301 => "001100100",
7302 => "001100101",
7303 => "001101011",
7304 => "001011111",
7305 => "001011100",
7306 => "001100001",
7307 => "001011111",
7308 => "001100011",
7309 => "001100010",
7310 => "001100101",
7311 => "001100000",
7312 => "001100110",
7313 => "001100100",
7314 => "001100110",
7315 => "001100111",
7316 => "001100101",
7317 => "001101100",
7318 => "001101101",
7319 => "001101100",
7320 => "001100111",
7321 => "001100110",
7322 => "001100011",
7323 => "000111101",
7324 => "001010011",
7325 => "001010100",
7326 => "001100111",
7327 => "001100011",
7328 => "001100111",
7329 => "011100010",
7330 => "011101110",
7331 => "011101111",
7332 => "001101110",
7333 => "001010100",
7334 => "001111011",
7335 => "010100000",
7336 => "010110100",
7337 => "010110111",
7338 => "010001111",
7339 => "010000010",
7340 => "010011011",
7341 => "010011011",
7342 => "010100011",
7343 => "011000100",
7344 => "010111101",
7345 => "010111101",
7346 => "011000110",
7347 => "011000100",
7348 => "011000001",
7349 => "011000001",
7350 => "011000101",
7351 => "011101011",
7352 => "011101011",
7353 => "011110110",
7354 => "011010011",
7355 => "011010000",
7356 => "011000010",
7357 => "011000011",
7358 => "011000101",
7359 => "010111111",
7360 => "010110010",
7361 => "010101111",
7362 => "010011110",
7363 => "010100000",
7364 => "010001100",
7365 => "010011101",
7366 => "010010101",
7367 => "010000010",
7368 => "001110111",
7369 => "001011110",
7370 => "001010011",
7371 => "001011101",
7372 => "001100101",
7373 => "001111110",
7374 => "011010100",
7375 => "011011000",
7376 => "011110100",
7377 => "011110011",
7378 => "011110100",
7379 => "011110011",
7380 => "011110100",
7381 => "011110011",
7382 => "011110100",
7383 => "011100101",
7384 => "011110000",
7385 => "011110010",
7386 => "011101110",
7387 => "011110011",
7388 => "011101110",
7389 => "011110101",
7390 => "011110100",
7391 => "011110010",
7392 => "011101110",
7393 => "011101110",
7394 => "011110011",
7395 => "011110000",
7396 => "011110000",
7397 => "011001010",
7398 => "001011100",
7399 => "001010111",
7400 => "001010100",
7401 => "001010010",
7402 => "001001110",
7403 => "001001111",
7404 => "001001010",
7405 => "001000001",
7406 => "010010011",
7407 => "011001000",
7408 => "011001101",
7409 => "011001011",
7410 => "011101110",
7411 => "011110000",
7412 => "010010010",
7413 => "001100001",
7414 => "001001010",
7415 => "001001011",
7416 => "001001111",
7417 => "001001100",
7418 => "001010001",
7419 => "001010001",
7420 => "001011100",
7421 => "001100000",
7422 => "001011011",
7423 => "001011101",
7424 => "001100110",
7425 => "001011111",
7426 => "001100010",
7427 => "001100001",
7428 => "001100000",
7429 => "001100001",
7430 => "001100000",
7431 => "001100101",
7432 => "001100010",
7433 => "001101010",
7434 => "001100110",
7435 => "001101000",
7436 => "001101011",
7437 => "001101111",
7438 => "001101110",
7439 => "001101101",
7440 => "001100001",
7441 => "001011101",
7442 => "001100011",
7443 => "001100001",
7444 => "001101001",
7445 => "001011110",
7446 => "001011111",
7447 => "001100100",
7448 => "001100001",
7449 => "001100111",
7450 => "001101100",
7451 => "001100001",
7452 => "001011111",
7453 => "001100010",
7454 => "001100101",
7455 => "001101011",
7456 => "001100110",
7457 => "011100100",
7458 => "010001000",
7459 => "010110010",
7460 => "001110010",
7461 => "001100110",
7462 => "001100100",
7463 => "001100101",
7464 => "001101001",
7465 => "001111110",
7466 => "010000011",
7467 => "001111001",
7468 => "010001011",
7469 => "010011000",
7470 => "010101000",
7471 => "010111101",
7472 => "011000100",
7473 => "011000000",
7474 => "011000011",
7475 => "011000010",
7476 => "011000010",
7477 => "010111101",
7478 => "010111111",
7479 => "011101101",
7480 => "011110010",
7481 => "011110101",
7482 => "011010100",
7483 => "011001010",
7484 => "011001010",
7485 => "011001110",
7486 => "010111110",
7487 => "010111011",
7488 => "011000001",
7489 => "011000100",
7490 => "011000001",
7491 => "010111111",
7492 => "001110111",
7493 => "000101111",
7494 => "010000010",
7495 => "010100000",
7496 => "010100000",
7497 => "010011101",
7498 => "010010111",
7499 => "010000110",
7500 => "001110101",
7501 => "010000111",
7502 => "011000011",
7503 => "011100011",
7504 => "011110010",
7505 => "011110000",
7506 => "011110100",
7507 => "011110110",
7508 => "011110100",
7509 => "011110000",
7510 => "011110100",
7511 => "011110110",
7512 => "011110101",
7513 => "011110000",
7514 => "011101111",
7515 => "011110011",
7516 => "011110100",
7517 => "011110011",
7518 => "011110011",
7519 => "011101111",
7520 => "011101111",
7521 => "011101011",
7522 => "011110100",
7523 => "011101111",
7524 => "011110001",
7525 => "011101010",
7526 => "001011001",
7527 => "001010101",
7528 => "001010101",
7529 => "001010001",
7530 => "001001111",
7531 => "001001011",
7532 => "001000101",
7533 => "001000011",
7534 => "010110101",
7535 => "011011011",
7536 => "011011001",
7537 => "011001100",
7538 => "010100000",
7539 => "010011011",
7540 => "010101100",
7541 => "001001011",
7542 => "001001001",
7543 => "001000110",
7544 => "001000110",
7545 => "001001011",
7546 => "001001001",
7547 => "001000001",
7548 => "001010011",
7549 => "010001001",
7550 => "001101001",
7551 => "001001101",
7552 => "001001011",
7553 => "001001111",
7554 => "001001011",
7555 => "001001111",
7556 => "001001011",
7557 => "001010000",
7558 => "001001110",
7559 => "001011000",
7560 => "001011101",
7561 => "001010111",
7562 => "001010111",
7563 => "001011110",
7564 => "001011011",
7565 => "001010011",
7566 => "001100000",
7567 => "001100010",
7568 => "001011011",
7569 => "001100011",
7570 => "001101001",
7571 => "001100111",
7572 => "001011100",
7573 => "001100111",
7574 => "001100101",
7575 => "001011010",
7576 => "001100100",
7577 => "001011111",
7578 => "001100101",
7579 => "001101011",
7580 => "001000101",
7581 => "001001000",
7582 => "001011101",
7583 => "001100111",
7584 => "001101010",
7585 => "010010011",
7586 => "001111010",
7587 => "010000000",
7588 => "001110010",
7589 => "001101001",
7590 => "001100110",
7591 => "001100101",
7592 => "001101000",
7593 => "001100111",
7594 => "010000101",
7595 => "010001000",
7596 => "001101111",
7597 => "001101100",
7598 => "001111010",
7599 => "010001011",
7600 => "010100101",
7601 => "010111001",
7602 => "011000000",
7603 => "010111011",
7604 => "011000001",
7605 => "011000011",
7606 => "010111111",
7607 => "011100000",
7608 => "011110001",
7609 => "011110010",
7610 => "011011000",
7611 => "011001101",
7612 => "011000111",
7613 => "011000111",
7614 => "011001001",
7615 => "011000111",
7616 => "010111110",
7617 => "011000110",
7618 => "011000001",
7619 => "010111110",
7620 => "010010011",
7621 => "000111100",
7622 => "010011110",
7623 => "011000000",
7624 => "010110110",
7625 => "010111000",
7626 => "010110101",
7627 => "010101000",
7628 => "010110101",
7629 => "010111001",
7630 => "011000000",
7631 => "011101100",
7632 => "011101110",
7633 => "011110010",
7634 => "011110110",
7635 => "011110111",
7636 => "011110110",
7637 => "011110110",
7638 => "011110101",
7639 => "011110011",
7640 => "011110110",
7641 => "011110011",
7642 => "011110000",
7643 => "011110011",
7644 => "011101111",
7645 => "011110001",
7646 => "011110100",
7647 => "011110001",
7648 => "011110010",
7649 => "011101111",
7650 => "011110101",
7651 => "011110011",
7652 => "011110101",
7653 => "011101011",
7654 => "001011101",
7655 => "001011000",
7656 => "001011000",
7657 => "001010011",
7658 => "001010100",
7659 => "001001101",
7660 => "001000100",
7661 => "001000011",
7662 => "001111000",
7663 => "010110110",
7664 => "010110000",
7665 => "010010001",
7666 => "010010011",
7667 => "010011001",
7668 => "010001110",
7669 => "001000101",
7670 => "001001101",
7671 => "001001110",
7672 => "001001110",
7673 => "001001001",
7674 => "001001110",
7675 => "001000100",
7676 => "001100000",
7677 => "010010001",
7678 => "001110100",
7679 => "001000110",
7680 => "001010001",
7681 => "001010001",
7682 => "001001100",
7683 => "001001001",
7684 => "001001101",
7685 => "001001001",
7686 => "001010011",
7687 => "001010010",
7688 => "001010010",
7689 => "001001100",
7690 => "001010000",
7691 => "001001111",
7692 => "001001110",
7693 => "001010011",
7694 => "001010011",
7695 => "001010111",
7696 => "001010110",
7697 => "001010011",
7698 => "001011011",
7699 => "001011110",
7700 => "001100011",
7701 => "001011011",
7702 => "001011111",
7703 => "001011101",
7704 => "001011010",
7705 => "001001111",
7706 => "001001111",
7707 => "001100011",
7708 => "001100010",
7709 => "001011100",
7710 => "001010011",
7711 => "001001101",
7712 => "001001010",
7713 => "010100110",
7714 => "010001000",
7715 => "010100001",
7716 => "001111010",
7717 => "001011111",
7718 => "001101010",
7719 => "001101001",
7720 => "001101101",
7721 => "001100110",
7722 => "010010000",
7723 => "010001110",
7724 => "001101011",
7725 => "001101000",
7726 => "001100111",
7727 => "001101010",
7728 => "001100110",
7729 => "001100001",
7730 => "001110000",
7731 => "010011001",
7732 => "010101001",
7733 => "010101110",
7734 => "010101101",
7735 => "011100001",
7736 => "011110001",
7737 => "011110000",
7738 => "011001111",
7739 => "011001110",
7740 => "011000101",
7741 => "011000011",
7742 => "011000111",
7743 => "011000010",
7744 => "011000001",
7745 => "011000001",
7746 => "011000011",
7747 => "011000101",
7748 => "010011110",
7749 => "000111110",
7750 => "010101111",
7751 => "011000111",
7752 => "011001001",
7753 => "010110001",
7754 => "010111111",
7755 => "011000001",
7756 => "011000000",
7757 => "011000001",
7758 => "011000001",
7759 => "011110011",
7760 => "011110111",
7761 => "011110100",
7762 => "011110011",
7763 => "011110100",
7764 => "011110111",
7765 => "011110100",
7766 => "011110100",
7767 => "011110110",
7768 => "011110011",
7769 => "011110010",
7770 => "011101000",
7771 => "011101011",
7772 => "011110100",
7773 => "011110011",
7774 => "011110011",
7775 => "011110001",
7776 => "011110011",
7777 => "011110011",
7778 => "011110100",
7779 => "011110100",
7780 => "011110011",
7781 => "011100111",
7782 => "001011000",
7783 => "001010100",
7784 => "001010011",
7785 => "001010101",
7786 => "010001111",
7787 => "010010100",
7788 => "001010100",
7789 => "001001010",
7790 => "001000001",
7791 => "010111001",
7792 => "011000011",
7793 => "001111101",
7794 => "010001110",
7795 => "010010011",
7796 => "001100110",
7797 => "001010110",
7798 => "001010101",
7799 => "001010100",
7800 => "001010111",
7801 => "001010011",
7802 => "001001100",
7803 => "001000101",
7804 => "001010001",
7805 => "010010001",
7806 => "001101001",
7807 => "001001011",
7808 => "001000111",
7809 => "001000101",
7810 => "000111111",
7811 => "001000001",
7812 => "000111110",
7813 => "000111100",
7814 => "001000010",
7815 => "000111110",
7816 => "001000101",
7817 => "001001111",
7818 => "001001010",
7819 => "001001110",
7820 => "001001100",
7821 => "001001100",
7822 => "001010000",
7823 => "001001111",
7824 => "001010010",
7825 => "001010100",
7826 => "001010001",
7827 => "001001100",
7828 => "001011101",
7829 => "001010000",
7830 => "001010101",
7831 => "001100001",
7832 => "001100000",
7833 => "001100011",
7834 => "001011100",
7835 => "001101000",
7836 => "001001000",
7837 => "001001101",
7838 => "001010101",
7839 => "001010110",
7840 => "001010110",
7841 => "001010000",
7842 => "001110010",
7843 => "010001001",
7844 => "010001101",
7845 => "001011111",
7846 => "001100001",
7847 => "001001001",
7848 => "001011010",
7849 => "001010111",
7850 => "001110100",
7851 => "001111000",
7852 => "001101101",
7853 => "001101101",
7854 => "001100111",
7855 => "001101101",
7856 => "001101011",
7857 => "001101010",
7858 => "001101100",
7859 => "001101000",
7860 => "001101000",
7861 => "001101011",
7862 => "001101001",
7863 => "001100110",
7864 => "001101100",
7865 => "010100000",
7866 => "010110010",
7867 => "010111010",
7868 => "011000101",
7869 => "011000111",
7870 => "011000011",
7871 => "010111100",
7872 => "010111110",
7873 => "010111010",
7874 => "011000011",
7875 => "010111110",
7876 => "010100110",
7877 => "001000110",
7878 => "010111000",
7879 => "010110001",
7880 => "010111101",
7881 => "011000110",
7882 => "010110101",
7883 => "010111101",
7884 => "010111110",
7885 => "010111100",
7886 => "011000000",
7887 => "011110100",
7888 => "011110100",
7889 => "011110100",
7890 => "011110101",
7891 => "011110111",
7892 => "011110011",
7893 => "011110101",
7894 => "011110011",
7895 => "011110101",
7896 => "011110010",
7897 => "011110110",
7898 => "011110100",
7899 => "011110000",
7900 => "011110010",
7901 => "011110010",
7902 => "011110100",
7903 => "011110010",
7904 => "011110010",
7905 => "011110011",
7906 => "011110100",
7907 => "011110011",
7908 => "011101111",
7909 => "011101100",
7910 => "001001111",
7911 => "001001110",
7912 => "001001111",
7913 => "001010001",
7914 => "010010101",
7915 => "010010011",
7916 => "001011100",
7917 => "001011101",
7918 => "001011110",
7919 => "010000001",
7920 => "010110001",
7921 => "001101111",
7922 => "010001010",
7923 => "010011001",
7924 => "001011111",
7925 => "001010111",
7926 => "001010100",
7927 => "001011100",
7928 => "001010110",
7929 => "001001100",
7930 => "001001001",
7931 => "001010000",
7932 => "001010010",
7933 => "001010101",
7934 => "001001101",
7935 => "001001001",
7936 => "001000011",
7937 => "000111011",
7938 => "001000000",
7939 => "000111100",
7940 => "000111110",
7941 => "001000001",
7942 => "000110111",
7943 => "000111001",
7944 => "000111101",
7945 => "001000101",
7946 => "001000110",
7947 => "001001101",
7948 => "001001110",
7949 => "001001011",
7950 => "001001010",
7951 => "001010111",
7952 => "001010100",
7953 => "001001101",
7954 => "001010011",
7955 => "001010011",
7956 => "001010101",
7957 => "001100010",
7958 => "001011100",
7959 => "001001110",
7960 => "001001011",
7961 => "001001101",
7962 => "001010001",
7963 => "001010111",
7964 => "001011010",
7965 => "001011111",
7966 => "001100000",
7967 => "001011110",
7968 => "001010110",
7969 => "001011000",
7970 => "001111010",
7971 => "010001111",
7972 => "010010011",
7973 => "001100100",
7974 => "001101001",
7975 => "001101001",
7976 => "001110010",
7977 => "001001101",
7978 => "001110110",
7979 => "001110111",
7980 => "001100000",
7981 => "001100000",
7982 => "001011110",
7983 => "001100100",
7984 => "001100100",
7985 => "001110100",
7986 => "001110001",
7987 => "001101011",
7988 => "001101010",
7989 => "001100111",
7990 => "001101100",
7991 => "001101000",
7992 => "001101001",
7993 => "001100111",
7994 => "001101011",
7995 => "001100111",
7996 => "001110001",
7997 => "010011110",
7998 => "010111001",
7999 => "011000001",
8000 => "011000100",
8001 => "011000001",
8002 => "010111101",
8003 => "011000010",
8004 => "011000000",
8005 => "011001001",
8006 => "010110100",
8007 => "011000011",
8008 => "011000000",
8009 => "010111111",
8010 => "011000100",
8011 => "010111101",
8012 => "010111100",
8013 => "011000001",
8014 => "011000100",
8015 => "011101010",
8016 => "011110001",
8017 => "011110101",
8018 => "011110001",
8019 => "011110110",
8020 => "011110101",
8021 => "011110010",
8022 => "011110100",
8023 => "011110101",
8024 => "011110010",
8025 => "011110101",
8026 => "011110011",
8027 => "011110010",
8028 => "011101101",
8029 => "011110010",
8030 => "011110000",
8031 => "011100110",
8032 => "011101110",
8033 => "011110000",
8034 => "011110001",
8035 => "011110000",
8036 => "011110000",
8037 => "011100011",
8038 => "001010110",
8039 => "001011110",
8040 => "001100000",
8041 => "001100101",
8042 => "010010101",
8043 => "010010010",
8044 => "001111100",
8045 => "001101001",
8046 => "001011101",
8047 => "001011011",
8048 => "001011011",
8049 => "001110000",
8050 => "010001011",
8051 => "010010011",
8052 => "001011110",
8053 => "001010110",
8054 => "001010111",
8055 => "001011001",
8056 => "001011000",
8057 => "001010001",
8058 => "001001111",
8059 => "001001100",
8060 => "001001010",
8061 => "001010010",
8062 => "001001101",
8063 => "001001101",
8064 => "001010101",
8065 => "001010011",
8066 => "001001111",
8067 => "001010011",
8068 => "001001100",
8069 => "001010001",
8070 => "001001011",
8071 => "001001011",
8072 => "001000111",
8073 => "001000101",
8074 => "001000111",
8075 => "001000101",
8076 => "000111111",
8077 => "000111100",
8078 => "000111110",
8079 => "001001010",
8080 => "001001011",
8081 => "001001010",
8082 => "001010000",
8083 => "001001101",
8084 => "001010011",
8085 => "001010101",
8086 => "001010110",
8087 => "001010010",
8088 => "001011011",
8089 => "001010111",
8090 => "001011000",
8091 => "001010001",
8092 => "001010101",
8093 => "001010100",
8094 => "001010000",
8095 => "001010101",
8096 => "001011010",
8097 => "001010110",
8098 => "001011001",
8099 => "001010110",
8100 => "001011101",
8101 => "001011010",
8102 => "001010101",
8103 => "001011110",
8104 => "001011111",
8105 => "001100001",
8106 => "001101001",
8107 => "001101101",
8108 => "001110000",
8109 => "001101101",
8110 => "001101110",
8111 => "001101100",
8112 => "001100001",
8113 => "001100010",
8114 => "001100100",
8115 => "001101001",
8116 => "001100010",
8117 => "001011111",
8118 => "001001010",
8119 => "001101001",
8120 => "001101101",
8121 => "001101111",
8122 => "001101111",
8123 => "001101101",
8124 => "001101110",
8125 => "001101011",
8126 => "001110000",
8127 => "001101100",
8128 => "010011001",
8129 => "010111001",
8130 => "011000000",
8131 => "011000011",
8132 => "010110111",
8133 => "011000101",
8134 => "011000110",
8135 => "011000011",
8136 => "011001100",
8137 => "011001100",
8138 => "011001101",
8139 => "011000101",
8140 => "010101010",
8141 => "011000001",
8142 => "010111011",
8143 => "011011010",
8144 => "011110000",
8145 => "011101111",
8146 => "011110001",
8147 => "011110010",
8148 => "011110011",
8149 => "011110101",
8150 => "011110100",
8151 => "011110001",
8152 => "011110000",
8153 => "011101111",
8154 => "011110010",
8155 => "011110011",
8156 => "011110100",
8157 => "011101111",
8158 => "011101110",
8159 => "011110101",
8160 => "011101000",
8161 => "011101111",
8162 => "011101110",
8163 => "011101111",
8164 => "011101110",
8165 => "011101000",
8166 => "001100100",
8167 => "001110110",
8168 => "001101101",
8169 => "000110011",
8170 => "010000111",
8171 => "010001011",
8172 => "010010011",
8173 => "010000100",
8174 => "001001101",
8175 => "000111110",
8176 => "000111110",
8177 => "001111101",
8178 => "010001111",
8179 => "010011001",
8180 => "001100110",
8181 => "001011000",
8182 => "001010100",
8183 => "001010001",
8184 => "001011000",
8185 => "001010011",
8186 => "001011011",
8187 => "001010100",
8188 => "001010100",
8189 => "001010001",
8190 => "001010100",
8191 => "001010000",
8192 => "001011010",
8193 => "001011000",
8194 => "001011001",
8195 => "001011000",
8196 => "001010111",
8197 => "001100000",
8198 => "001011000",
8199 => "001011000",
8200 => "001011000",
8201 => "001010101",
8202 => "001010010",
8203 => "001010010",
8204 => "001011000",
8205 => "001010110",
8206 => "001010010",
8207 => "001001111",
8208 => "001001000",
8209 => "001001001",
8210 => "001001101",
8211 => "001001111",
8212 => "001010011",
8213 => "001001100",
8214 => "001010000",
8215 => "001010001",
8216 => "001010000",
8217 => "001001011",
8218 => "001001011",
8219 => "001000101",
8220 => "001001110",
8221 => "001000111",
8222 => "001001011",
8223 => "001001001",
8224 => "001001111",
8225 => "001010000",
8226 => "001011011",
8227 => "001011000",
8228 => "001010111",
8229 => "001011000",
8230 => "001010001",
8231 => "001010011",
8232 => "001010110",
8233 => "001011000",
8234 => "001001010",
8235 => "001000111",
8236 => "001011000",
8237 => "001010101",
8238 => "001011011",
8239 => "001100101",
8240 => "001101010",
8241 => "001100111",
8242 => "001101011",
8243 => "001101001",
8244 => "001101010",
8245 => "001100111",
8246 => "001111000",
8247 => "001100001",
8248 => "001100100",
8249 => "001100000",
8250 => "001100110",
8251 => "001101011",
8252 => "001110111",
8253 => "001101000",
8254 => "001101001",
8255 => "001101011",
8256 => "001110100",
8257 => "001110101",
8258 => "001111001",
8259 => "010000100",
8260 => "010101011",
8261 => "011000001",
8262 => "010111001",
8263 => "010111100",
8264 => "011001001",
8265 => "010110001",
8266 => "011001000",
8267 => "011001001",
8268 => "010010001",
8269 => "010011110",
8270 => "010111110",
8271 => "011101110",
8272 => "011101101",
8273 => "011110010",
8274 => "011110010",
8275 => "011110011",
8276 => "011110010",
8277 => "011110010",
8278 => "011101101",
8279 => "011110010",
8280 => "011110011",
8281 => "011101101",
8282 => "011101110",
8283 => "011101111",
8284 => "011110100",
8285 => "011110010",
8286 => "011110001",
8287 => "011110011",
8288 => "011101110",
8289 => "011101010",
8290 => "011110001",
8291 => "011101000",
8292 => "011101011",
8293 => "011110001",
8294 => "001011111",
8295 => "001111100",
8296 => "010000001",
8297 => "001011011",
8298 => "001011101",
8299 => "010001001",
8300 => "010011011",
8301 => "010000101",
8302 => "001100000",
8303 => "001010110",
8304 => "001001110",
8305 => "001011110",
8306 => "001100110",
8307 => "001011010",
8308 => "001010111",
8309 => "001011010",
8310 => "001011001",
8311 => "001011100",
8312 => "001010101",
8313 => "001010110",
8314 => "001011011",
8315 => "001010111",
8316 => "001010011",
8317 => "001010100",
8318 => "001010010",
8319 => "001010011",
8320 => "001010100",
8321 => "001011000",
8322 => "001011100",
8323 => "001010101",
8324 => "001100001",
8325 => "001011100",
8326 => "001011101",
8327 => "001011100",
8328 => "001011011",
8329 => "001011011",
8330 => "001100000",
8331 => "001011111",
8332 => "001011110",
8333 => "001011000",
8334 => "001010110",
8335 => "001011101",
8336 => "001010100",
8337 => "001010101",
8338 => "001011011",
8339 => "001010110",
8340 => "001010100",
8341 => "001010101",
8342 => "001001100",
8343 => "001001000",
8344 => "001001100",
8345 => "001010100",
8346 => "001001100",
8347 => "001001110",
8348 => "001001000",
8349 => "001001100",
8350 => "001000011",
8351 => "001000111",
8352 => "001001011",
8353 => "001000000",
8354 => "001010100",
8355 => "001001111",
8356 => "001001101",
8357 => "001010110",
8358 => "001001101",
8359 => "001001101",
8360 => "001010011",
8361 => "001011000",
8362 => "001010011",
8363 => "001001110",
8364 => "001011000",
8365 => "001011001",
8366 => "001010100",
8367 => "001011110",
8368 => "001100000",
8369 => "001011110",
8370 => "001011111",
8371 => "001011111",
8372 => "001100110",
8373 => "001100100",
8374 => "001010001",
8375 => "001100001",
8376 => "001100011",
8377 => "001011011",
8378 => "001100001",
8379 => "001100001",
8380 => "001101000",
8381 => "001100010",
8382 => "001110101",
8383 => "001100100",
8384 => "001101001",
8385 => "001100111",
8386 => "001101111",
8387 => "001100011",
8388 => "001100111",
8389 => "001101111",
8390 => "010000000",
8391 => "010011000",
8392 => "010011001",
8393 => "010100010",
8394 => "010100111",
8395 => "010101101",
8396 => "010000101",
8397 => "010011011",
8398 => "010101100",
8399 => "011101011",
8400 => "011110000",
8401 => "011110100",
8402 => "011110000",
8403 => "011101101",
8404 => "011101111",
8405 => "011110010",
8406 => "011110011",
8407 => "011110100",
8408 => "011110100",
8409 => "011101100",
8410 => "011110000",
8411 => "011110101",
8412 => "011011001",
8413 => "010111010",
8414 => "010111100",
8415 => "011110010",
8416 => "011110001",
8417 => "011110101",
8418 => "010111111",
8419 => "010111110",
8420 => "011100110",
8421 => "011101011",
8422 => "001110001",
8423 => "001111111",
8424 => "010000001",
8425 => "001011010",
8426 => "001100100",
8427 => "010001110",
8428 => "010011101",
8429 => "010000011",
8430 => "001100000",
8431 => "001011110",
8432 => "001011000",
8433 => "001010101",
8434 => "001011001",
8435 => "001011001",
8436 => "001010010",
8437 => "010000101",
8438 => "001100111",
8439 => "001011110",
8440 => "001100001",
8441 => "001011111",
8442 => "001011100",
8443 => "001011001",
8444 => "001010101",
8445 => "001010101",
8446 => "001010101",
8447 => "001011000",
8448 => "001011010",
8449 => "001011110",
8450 => "001011110",
8451 => "001010110",
8452 => "001010101",
8453 => "001011100",
8454 => "001010011",
8455 => "001010101",
8456 => "001011011",
8457 => "001010111",
8458 => "001010110",
8459 => "001011101",
8460 => "001011111",
8461 => "001011110",
8462 => "001011101",
8463 => "001011101",
8464 => "001011111",
8465 => "001011100",
8466 => "001011110",
8467 => "001011111",
8468 => "001011111",
8469 => "001011010",
8470 => "001011010",
8471 => "001010100",
8472 => "001010010",
8473 => "001010101",
8474 => "001010010",
8475 => "001010101",
8476 => "001001000",
8477 => "001001011",
8478 => "001001011",
8479 => "001001101",
8480 => "001001100",
8481 => "000111101",
8482 => "001000011",
8483 => "001000100",
8484 => "001001011",
8485 => "001000110",
8486 => "001000010",
8487 => "001000101",
8488 => "001000100",
8489 => "001001000",
8490 => "001000101",
8491 => "001010110",
8492 => "001010100",
8493 => "001010101",
8494 => "001010001",
8495 => "001010011",
8496 => "001010101",
8497 => "001100001",
8498 => "001010001",
8499 => "001001101",
8500 => "001010000",
8501 => "001010001",
8502 => "001011011",
8503 => "001011011",
8504 => "001001110",
8505 => "001010011",
8506 => "001100100",
8507 => "001100001",
8508 => "001011111",
8509 => "001011001",
8510 => "001011100",
8511 => "001100110",
8512 => "001101011",
8513 => "001100100",
8514 => "001101000",
8515 => "001101000",
8516 => "001100001",
8517 => "001100010",
8518 => "001110100",
8519 => "010001010",
8520 => "001111011",
8521 => "001010100",
8522 => "000111110",
8523 => "000111011",
8524 => "001111011",
8525 => "010010110",
8526 => "001111011",
8527 => "010011111",
8528 => "011000010",
8529 => "010110011",
8530 => "010011001",
8531 => "010011111",
8532 => "011000001",
8533 => "011100000",
8534 => "011111100",
8535 => "011111000",
8536 => "011110101",
8537 => "011110111",
8538 => "011110110",
8539 => "011011101",
8540 => "010101010",
8541 => "010110101",
8542 => "010111101",
8543 => "010001101",
8544 => "010000011",
8545 => "001110000",
8546 => "001111011",
8547 => "001111011",
8548 => "001101000",
8549 => "001100101",
8550 => "001100011",
8551 => "001111101",
8552 => "010000110",
8553 => "010000000",
8554 => "001101110",
8555 => "010001111",
8556 => "010011100",
8557 => "010000011",
8558 => "001100001",
8559 => "001011100",
8560 => "001100000",
8561 => "001011111",
8562 => "001110100",
8563 => "001101110",
8564 => "001101110",
8565 => "010001000",
8566 => "001111001",
8567 => "001011011",
8568 => "001011010",
8569 => "001010111",
8570 => "001011010",
8571 => "001011100",
8572 => "001011101",
8573 => "001011010",
8574 => "001011010",
8575 => "001011000",
8576 => "001010101",
8577 => "001010110",
8578 => "001011011",
8579 => "001010101",
8580 => "001011101",
8581 => "001011000",
8582 => "001011001",
8583 => "001011011",
8584 => "001011011",
8585 => "001010010",
8586 => "001100000",
8587 => "001010110",
8588 => "001010011",
8589 => "001011110",
8590 => "001011110",
8591 => "001011001",
8592 => "001011100",
8593 => "001011110",
8594 => "001011110",
8595 => "001011111",
8596 => "001011101",
8597 => "001011100",
8598 => "001011100",
8599 => "001011001",
8600 => "001010000",
8601 => "001011100",
8602 => "001011010",
8603 => "001011001",
8604 => "001011100",
8605 => "001010111",
8606 => "001010011",
8607 => "001001011",
8608 => "001001001",
8609 => "001001101",
8610 => "001001011",
8611 => "001001100",
8612 => "001001111",
8613 => "001001100",
8614 => "001000010",
8615 => "001000110",
8616 => "001001000",
8617 => "001000001",
8618 => "000110011",
8619 => "000111000",
8620 => "001000110",
8621 => "001001000",
8622 => "001000000",
8623 => "001000100",
8624 => "001001000",
8625 => "001001000",
8626 => "001001001",
8627 => "001001111",
8628 => "001010111",
8629 => "001011000",
8630 => "001010010",
8631 => "001010001",
8632 => "001011011",
8633 => "001010111",
8634 => "001001001",
8635 => "001000011",
8636 => "001001010",
8637 => "001100000",
8638 => "001101110",
8639 => "001100010",
8640 => "001100100",
8641 => "001011011",
8642 => "001011010",
8643 => "001010000",
8644 => "001011110",
8645 => "001011010",
8646 => "001011110",
8647 => "001110010",
8648 => "001101000",
8649 => "001101110",
8650 => "001011110",
8651 => "001001000",
8652 => "001101011",
8653 => "010001111",
8654 => "010000111",
8655 => "001111000",
8656 => "001111000",
8657 => "010001001",
8658 => "010011111",
8659 => "010001111",
8660 => "010000110",
8661 => "001110011",
8662 => "001101100",
8663 => "001111111",
8664 => "010001000",
8665 => "001111001",
8666 => "001110111",
8667 => "001100111",
8668 => "001111111",
8669 => "010111001",
8670 => "010111100",
8671 => "001100100",
8672 => "001100110",
8673 => "001101001",
8674 => "001110111",
8675 => "001110101",
8676 => "001100101",
8677 => "001100101",
8678 => "001101000",
8679 => "001111001",
8680 => "001111111",
8681 => "010010001",
8682 => "001100011",
8683 => "010010000",
8684 => "010011101",
8685 => "001111011",
8686 => "001011111",
8687 => "001100010",
8688 => "001100100",
8689 => "001100001",
8690 => "001111000",
8691 => "001111000",
8692 => "001100001",
8693 => "001100111",
8694 => "001011010",
8695 => "001011001",
8696 => "001100010",
8697 => "001100001",
8698 => "001011101",
8699 => "001011010",
8700 => "001011101",
8701 => "001011011",
8702 => "001010101",
8703 => "001011001",
8704 => "001011000",
8705 => "001011001",
8706 => "001011010",
8707 => "001010111",
8708 => "001010010",
8709 => "001010111",
8710 => "001011011",
8711 => "001100000",
8712 => "001010111",
8713 => "001011010",
8714 => "001011010",
8715 => "001010010",
8716 => "001011010",
8717 => "001010001",
8718 => "001001101",
8719 => "001010010",
8720 => "001011000",
8721 => "001011111",
8722 => "001011001",
8723 => "001010111",
8724 => "001011100",
8725 => "001100000",
8726 => "001011111",
8727 => "001100001",
8728 => "001100000",
8729 => "001011111",
8730 => "001100001",
8731 => "001100001",
8732 => "001011111",
8733 => "001011110",
8734 => "001100001",
8735 => "001100001",
8736 => "001011110",
8737 => "001011100",
8738 => "001100110",
8739 => "001011100",
8740 => "001011001",
8741 => "001010000",
8742 => "001001101",
8743 => "001001101",
8744 => "001010000",
8745 => "001010101",
8746 => "001001101",
8747 => "001000010",
8748 => "001000100",
8749 => "001000011",
8750 => "001000101",
8751 => "001001100",
8752 => "001001101",
8753 => "001001001",
8754 => "001001111",
8755 => "000111110",
8756 => "001000001",
8757 => "001000100",
8758 => "001011000",
8759 => "001010111",
8760 => "001010101",
8761 => "001101100",
8762 => "001110100",
8763 => "001011100",
8764 => "001001001",
8765 => "001101111",
8766 => "010000111",
8767 => "001011100",
8768 => "001001010",
8769 => "001011111",
8770 => "001010111",
8771 => "001011110",
8772 => "001011000",
8773 => "001011000",
8774 => "001010111",
8775 => "001010100",
8776 => "001011010",
8777 => "001011010",
8778 => "001011101",
8779 => "001011011",
8780 => "001010110",
8781 => "001011000",
8782 => "001011010",
8783 => "001100110",
8784 => "001100010",
8785 => "001101100",
8786 => "001101011",
8787 => "001101111",
8788 => "001100111",
8789 => "001101011",
8790 => "001101001",
8791 => "001101001",
8792 => "001101010",
8793 => "001100110",
8794 => "001101001",
8795 => "001101101",
8796 => "001111111",
8797 => "010011110",
8798 => "010100101",
8799 => "001100110",
8800 => "001100010",
8801 => "001101011",
8802 => "001111000",
8803 => "001110011",
8804 => "001011101",
8805 => "001011111",
8806 => "001101111",
8807 => "001111000",
8808 => "010000001",
8809 => "010010000",
8810 => "001101011",
8811 => "010010010",
8812 => "010011001",
8813 => "001111011",
8814 => "001011101",
8815 => "001011101",
8816 => "001011110",
8817 => "001101011",
8818 => "001111010",
8819 => "001110000",
8820 => "001011111",
8821 => "001010111",
8822 => "001011111",
8823 => "001010111",
8824 => "001011100",
8825 => "001011011",
8826 => "001011110",
8827 => "001011001",
8828 => "001011100",
8829 => "001011010",
8830 => "001011010",
8831 => "001011011",
8832 => "001100011",
8833 => "001100000",
8834 => "001011111",
8835 => "001010111",
8836 => "001011100",
8837 => "001011011",
8838 => "001010000",
8839 => "001010101",
8840 => "001100000",
8841 => "001100001",
8842 => "001011001",
8843 => "001011100",
8844 => "001010100",
8845 => "001010111",
8846 => "001010101",
8847 => "001010110",
8848 => "001011101",
8849 => "001011101",
8850 => "001011011",
8851 => "001011101",
8852 => "001011000",
8853 => "001010101",
8854 => "001100011",
8855 => "001010011",
8856 => "001011101",
8857 => "001011110",
8858 => "001100001",
8859 => "001100010",
8860 => "001011111",
8861 => "001100000",
8862 => "001011111",
8863 => "001011110",
8864 => "001011111",
8865 => "001011100",
8866 => "001011100",
8867 => "001011110",
8868 => "001011000",
8869 => "001011001",
8870 => "001011110",
8871 => "001011100",
8872 => "001010010",
8873 => "001010101",
8874 => "001010001",
8875 => "001010101",
8876 => "001010001",
8877 => "001001010",
8878 => "001010101",
8879 => "001010001",
8880 => "001010111",
8881 => "001010111",
8882 => "001001101",
8883 => "001001101",
8884 => "001000111",
8885 => "001000001",
8886 => "001000011",
8887 => "001000011",
8888 => "000111101",
8889 => "001001101",
8890 => "001011000",
8891 => "001101111",
8892 => "001110010",
8893 => "001010011",
8894 => "001110110",
8895 => "001100011",
8896 => "001011000",
8897 => "001001101",
8898 => "001001101",
8899 => "001001001",
8900 => "001011010",
8901 => "001100010",
8902 => "001110101",
8903 => "001100111",
8904 => "001010110",
8905 => "001010110",
8906 => "001010100",
8907 => "001010101",
8908 => "001011001",
8909 => "001100001",
8910 => "001100100",
8911 => "001101000",
8912 => "001100100",
8913 => "001100000",
8914 => "001011110",
8915 => "001100000",
8916 => "001011111",
8917 => "001100000",
8918 => "001100110",
8919 => "001101110",
8920 => "001100111",
8921 => "001101001",
8922 => "001101011",
8923 => "001100100",
8924 => "001011110",
8925 => "001011010",
8926 => "001011101",
8927 => "001100101",
8928 => "001100011",
8929 => "001100101",
8930 => "001101100",
8931 => "001101111",
8932 => "001100001",
8933 => "001100100",
8934 => "001100011",
8935 => "001101000",
8936 => "010000101",
8937 => "010001110",
8938 => "001100001",
8939 => "001011101",
8940 => "001011000",
8941 => "001011010",
8942 => "001011111",
8943 => "001011110",
8944 => "001001111",
8945 => "001011011",
8946 => "001010100",
8947 => "001011111",
8948 => "001011101",
8949 => "001010111",
8950 => "001010101",
8951 => "001011101",
8952 => "001011101",
8953 => "001011100",
8954 => "001011010",
8955 => "001011110",
8956 => "001011100",
8957 => "001011101",
8958 => "001010110",
8959 => "001100100",
8960 => "001100011",
8961 => "001100001",
8962 => "001100100",
8963 => "001100001",
8964 => "001010011",
8965 => "001011000",
8966 => "001010111",
8967 => "001011110",
8968 => "001011101",
8969 => "001100001",
8970 => "001011100",
8971 => "001011000",
8972 => "001001110",
8973 => "001001110",
8974 => "001010010",
8975 => "001100100",
8976 => "001101101",
8977 => "001011101",
8978 => "001011111",
8979 => "001011101",
8980 => "001010011",
8981 => "001011011",
8982 => "001011011",
8983 => "001100111",
8984 => "001100010",
8985 => "001100000",
8986 => "001100001",
8987 => "001011110",
8988 => "001011011",
8989 => "001100000",
8990 => "001011001",
8991 => "001100001",
8992 => "001011111",
8993 => "001100011",
8994 => "001100011",
8995 => "001100011",
8996 => "001100011",
8997 => "001100010",
8998 => "001011111",
8999 => "001011110",
9000 => "001011101",
9001 => "001011010",
9002 => "001100000",
9003 => "001011100",
9004 => "001011110",
9005 => "001011000",
9006 => "001011000",
9007 => "001100000",
9008 => "001011100",
9009 => "001010101",
9010 => "001010010",
9011 => "001001111",
9012 => "001001110",
9013 => "001000111",
9014 => "001000000",
9015 => "001001001",
9016 => "001001000",
9017 => "001001000",
9018 => "001001111",
9019 => "001000011",
9020 => "001001110",
9021 => "001001010",
9022 => "001001101",
9023 => "001011101",
9024 => "001110001",
9025 => "001110011",
9026 => "001011110",
9027 => "001100100",
9028 => "001011100",
9029 => "001001010",
9030 => "001001100",
9031 => "001000110",
9032 => "001001001",
9033 => "001000001",
9034 => "001000011",
9035 => "001010101",
9036 => "001011111",
9037 => "001011100",
9038 => "001010101",
9039 => "001011000",
9040 => "001011011",
9041 => "001011111",
9042 => "001011011",
9043 => "001011100",
9044 => "001011110",
9045 => "001011110",
9046 => "001011100",
9047 => "001011010",
9048 => "001010111",
9049 => "001100111",
9050 => "001100000",
9051 => "001100010",
9052 => "001100011",
9053 => "001100100",
9054 => "001100001",
9055 => "001100011",
9056 => "001100100",
9057 => "001100001",
9058 => "001100001",
9059 => "001011111",
9060 => "001011111",
9061 => "001100100",
9062 => "001011100",
9063 => "001011110",
9064 => "001110111",
9065 => "001111100",
9066 => "001101010",
9067 => "001100010",
9068 => "001011110",
9069 => "001011100",
9070 => "001100010",
9071 => "001100110",
9072 => "001100000",
9073 => "001011111",
9074 => "001100010",
9075 => "001011111",
9076 => "001100000",
9077 => "001100001",
9078 => "001011011",
9079 => "001011111",
9080 => "001011100",
9081 => "001010110",
9082 => "001011100",
9083 => "001010101",
9084 => "001010110",
9085 => "001011000",
9086 => "001010111",
9087 => "001011001",
9088 => "001101000",
9089 => "001100010",
9090 => "001100111",
9091 => "001100100",
9092 => "001100001",
9093 => "001100001",
9094 => "001101001",
9095 => "001100000",
9096 => "001100010",
9097 => "001100010",
9098 => "001101010",
9099 => "001100111",
9100 => "001100001",
9101 => "001011000",
9102 => "001011000",
9103 => "001010110",
9104 => "001011000",
9105 => "001010010",
9106 => "001011011",
9107 => "001100110",
9108 => "001011010",
9109 => "001011010",
9110 => "001011001",
9111 => "001101000",
9112 => "001011011",
9113 => "001011000",
9114 => "001011100",
9115 => "001100000",
9116 => "001100110",
9117 => "001100011",
9118 => "001100100",
9119 => "001100000",
9120 => "001100011",
9121 => "001100010",
9122 => "001011111",
9123 => "001011111",
9124 => "001011110",
9125 => "001001100",
9126 => "001001111",
9127 => "001100001",
9128 => "001101010",
9129 => "001100110",
9130 => "001100001",
9131 => "001011100",
9132 => "001100000",
9133 => "001011110",
9134 => "001011100",
9135 => "001011001",
9136 => "001010110",
9137 => "001100001",
9138 => "001011110",
9139 => "001011011",
9140 => "001011100",
9141 => "001011010",
9142 => "001011000",
9143 => "001011000",
9144 => "001010010",
9145 => "001001001",
9146 => "001001000",
9147 => "001010001",
9148 => "001001001",
9149 => "001001101",
9150 => "001001011",
9151 => "001000100",
9152 => "001001111",
9153 => "001010100",
9154 => "001010011",
9155 => "001010110",
9156 => "001001011",
9157 => "001010001",
9158 => "001011001",
9159 => "001010101",
9160 => "001010011",
9161 => "001011100",
9162 => "001001110",
9163 => "001000010",
9164 => "001010100",
9165 => "001010010",
9166 => "001001001",
9167 => "001010100",
9168 => "001010010",
9169 => "001011000",
9170 => "001011010",
9171 => "001011111",
9172 => "001011010",
9173 => "001010111",
9174 => "001010101",
9175 => "001010010",
9176 => "001010001",
9177 => "001001111",
9178 => "001010111",
9179 => "001011001",
9180 => "001011100",
9181 => "001100110",
9182 => "001100110",
9183 => "001100100",
9184 => "001100000",
9185 => "001011111",
9186 => "001011010",
9187 => "001011111",
9188 => "001100000",
9189 => "001100110",
9190 => "001100000",
9191 => "001011101",
9192 => "001100010",
9193 => "001011110",
9194 => "001011010",
9195 => "001011011",
9196 => "001011100",
9197 => "001011100",
9198 => "001100100",
9199 => "001011010",
9200 => "001100011",
9201 => "001011001",
9202 => "001011001",
9203 => "001011110",
9204 => "001011010",
9205 => "001011101",
9206 => "001010110",
9207 => "001011110",
9208 => "001010100",
9209 => "001010100",
9210 => "001001001",
9211 => "001001111",
9212 => "001011000",
9213 => "001010000",
9214 => "001010110",
9215 => "001011000",
9216 => "001101011",
9217 => "010001001",
9218 => "001101001",
9219 => "001110101",
9220 => "010000111",
9221 => "010010110",
9222 => "010001100",
9223 => "010011110",
9224 => "001111000",
9225 => "001001110",
9226 => "001101000",
9227 => "001101000",
9228 => "001100011",
9229 => "001100110",
9230 => "001100001",
9231 => "001101001",
9232 => "001011101",
9233 => "001100010",
9234 => "001011111",
9235 => "001011011",
9236 => "001011110",
9237 => "001100111",
9238 => "001100110",
9239 => "001011110",
9240 => "001011101",
9241 => "001100001",
9242 => "001100011",
9243 => "001100001",
9244 => "001100011",
9245 => "001011000",
9246 => "001100000",
9247 => "001011010",
9248 => "001011001",
9249 => "001100001",
9250 => "001100011",
9251 => "001100010",
9252 => "001100011",
9253 => "001100101",
9254 => "001100100",
9255 => "001100001",
9256 => "001100010",
9257 => "001100101",
9258 => "001100000",
9259 => "001100011",
9260 => "001100101",
9261 => "001100010",
9262 => "001100111",
9263 => "001100101",
9264 => "001100011",
9265 => "001100101",
9266 => "001100100",
9267 => "001100100",
9268 => "001011101",
9269 => "001011111",
9270 => "001011010",
9271 => "001001111",
9272 => "001010000",
9273 => "001010001",
9274 => "001100000",
9275 => "001011000",
9276 => "001010000",
9277 => "001001111",
9278 => "001010100",
9279 => "001010111",
9280 => "001010001",
9281 => "001001111",
9282 => "001011011",
9283 => "001010011",
9284 => "001001100",
9285 => "001010100",
9286 => "001010101",
9287 => "001000001",
9288 => "000110010",
9289 => "000111011",
9290 => "001000010",
9291 => "000111101",
9292 => "001000010",
9293 => "001000110",
9294 => "001001001",
9295 => "001001100",
9296 => "001001100",
9297 => "001001100",
9298 => "001010000",
9299 => "001010111",
9300 => "001010011",
9301 => "001011010",
9302 => "000111101",
9303 => "001000111",
9304 => "001010101",
9305 => "001010011",
9306 => "001010011",
9307 => "001010010",
9308 => "001101010",
9309 => "001011100",
9310 => "001010111",
9311 => "001011110",
9312 => "001100101",
9313 => "001010111",
9314 => "001001101",
9315 => "001010000",
9316 => "001011010",
9317 => "001101001",
9318 => "001101011",
9319 => "001011111",
9320 => "001011101",
9321 => "001100000",
9322 => "001011101",
9323 => "001011110",
9324 => "001011111",
9325 => "001100001",
9326 => "001100000",
9327 => "001011111",
9328 => "001100101",
9329 => "001011100",
9330 => "001101010",
9331 => "001011100",
9332 => "001010101",
9333 => "001011101",
9334 => "001011101",
9335 => "001011100",
9336 => "001010000",
9337 => "001100000",
9338 => "001010111",
9339 => "001011110",
9340 => "001011100",
9341 => "001010011",
9342 => "001001100",
9343 => "001001100",
9344 => "001101011",
9345 => "001011000",
9346 => "001101100",
9347 => "001010110",
9348 => "001001000",
9349 => "001010101",
9350 => "000111100",
9351 => "001101110",
9352 => "001110111",
9353 => "000111111",
9354 => "001010001",
9355 => "001100010",
9356 => "001101101",
9357 => "001100100",
9358 => "001100000",
9359 => "001100001",
9360 => "001011011",
9361 => "001100111",
9362 => "001100011",
9363 => "001101001",
9364 => "001100101",
9365 => "001101011",
9366 => "001100111",
9367 => "001100110",
9368 => "001100011",
9369 => "001011101",
9370 => "001011010",
9371 => "001100111",
9372 => "001100101",
9373 => "001100011",
9374 => "001100011",
9375 => "001100110",
9376 => "001011111",
9377 => "001100010",
9378 => "001010010",
9379 => "001011110",
9380 => "001101001",
9381 => "001100110",
9382 => "001100010",
9383 => "001100000",
9384 => "001101000",
9385 => "001101010",
9386 => "001100100",
9387 => "001100001",
9388 => "001100011",
9389 => "001011010",
9390 => "001100001",
9391 => "001011011",
9392 => "001011111",
9393 => "001100010",
9394 => "001100110",
9395 => "001101001",
9396 => "001101011",
9397 => "001101000",
9398 => "001100011",
9399 => "001100000",
9400 => "001100010",
9401 => "001011111",
9402 => "001011101",
9403 => "001011111",
9404 => "001011010",
9405 => "001011101",
9406 => "001100000",
9407 => "001011110",
9408 => "001010111",
9409 => "001011000",
9410 => "001011010",
9411 => "001010110",
9412 => "001010011",
9413 => "001010001",
9414 => "001001100",
9415 => "001001001",
9416 => "001001000",
9417 => "001000010",
9418 => "000111110",
9419 => "001000000",
9420 => "001000011",
9421 => "001000111",
9422 => "001001100",
9423 => "001010001",
9424 => "001000011",
9425 => "001000010",
9426 => "001000010",
9427 => "001000100",
9428 => "001000011",
9429 => "001001111",
9430 => "001001101",
9431 => "001001111",
9432 => "001011110",
9433 => "001001010",
9434 => "001010011",
9435 => "001001011",
9436 => "001101001",
9437 => "001011110",
9438 => "001100000",
9439 => "001011110",
9440 => "001011011",
9441 => "001100010",
9442 => "001011010",
9443 => "001000101",
9444 => "001100011",
9445 => "001100111",
9446 => "001101010",
9447 => "001100100",
9448 => "001100001",
9449 => "001011010",
9450 => "001011001",
9451 => "001011111",
9452 => "001011001",
9453 => "001100100",
9454 => "001100011",
9455 => "001010111",
9456 => "001100010",
9457 => "001011100",
9458 => "001110000",
9459 => "001100001",
9460 => "001100001",
9461 => "001011001",
9462 => "001011100",
9463 => "001011111",
9464 => "001001111",
9465 => "001011110",
9466 => "001011000",
9467 => "001010011",
9468 => "001001011",
9469 => "001001111",
9470 => "001001101",
9471 => "001001111",
9472 => "001010010",
9473 => "001110001",
9474 => "001010110",
9475 => "001010010",
9476 => "001000100",
9477 => "001001000",
9478 => "001001001",
9479 => "001001011",
9480 => "001010001",
9481 => "001010001",
9482 => "001000000",
9483 => "001010111",
9484 => "001110001",
9485 => "001100110",
9486 => "001100101",
9487 => "001110011",
9488 => "001110000",
9489 => "001101111",
9490 => "001100010",
9491 => "001100011",
9492 => "001100101",
9493 => "001101001",
9494 => "001101110",
9495 => "001100011",
9496 => "001011100",
9497 => "001101000",
9498 => "001011110",
9499 => "001011000",
9500 => "001011011",
9501 => "001011011",
9502 => "001010111",
9503 => "001011101",
9504 => "001011100",
9505 => "001010110",
9506 => "001100111",
9507 => "001100110",
9508 => "001100011",
9509 => "001011100",
9510 => "001011111",
9511 => "001100010",
9512 => "001101101",
9513 => "001101000",
9514 => "001011001",
9515 => "001100011",
9516 => "001100101",
9517 => "001011101",
9518 => "001100100",
9519 => "001010011",
9520 => "001011100",
9521 => "001100010",
9522 => "001100011",
9523 => "001011110",
9524 => "001010110",
9525 => "001010001",
9526 => "001011101",
9527 => "001100001",
9528 => "001011011",
9529 => "001100101",
9530 => "001100001",
9531 => "001100000",
9532 => "001100000",
9533 => "001100100",
9534 => "001100000",
9535 => "001100001",
9536 => "001100011",
9537 => "001100100",
9538 => "001011111",
9539 => "001011110",
9540 => "001011110",
9541 => "001011010",
9542 => "001010111",
9543 => "001010000",
9544 => "001001010",
9545 => "001001011",
9546 => "001010111",
9547 => "001000111",
9548 => "001000111",
9549 => "001010100",
9550 => "001001001",
9551 => "001001000",
9552 => "000111110",
9553 => "001000101",
9554 => "001000111",
9555 => "001000110",
9556 => "001001011",
9557 => "001001110",
9558 => "001001011",
9559 => "001010101",
9560 => "001001100",
9561 => "001000111",
9562 => "001010101",
9563 => "001011001",
9564 => "001100010",
9565 => "001100001",
9566 => "001100100",
9567 => "001011010",
9568 => "001011110",
9569 => "001011110",
9570 => "001010111",
9571 => "001011111",
9572 => "001100110",
9573 => "001101000",
9574 => "001011010",
9575 => "001101101",
9576 => "001111000",
9577 => "001101100",
9578 => "001111001",
9579 => "001011000",
9580 => "001011010",
9581 => "001100011",
9582 => "001011111",
9583 => "001011000",
9584 => "001011100",
9585 => "001010100",
9586 => "001010001",
9587 => "001010010",
9588 => "001011011",
9589 => "001011001",
9590 => "001010101",
9591 => "001010110",
9592 => "001010100",
9593 => "001010101",
9594 => "001010000",
9595 => "001001111",
9596 => "001001011",
9597 => "001010101",
9598 => "001010011",
9599 => "001000110",
9600 => "001110111",
9601 => "001001100",
9602 => "000110110",
9603 => "000100101",
9604 => "001001111",
9605 => "000111111",
9606 => "001010000",
9607 => "001011111",
9608 => "001000101",
9609 => "001001100",
9610 => "001001100",
9611 => "001001000",
9612 => "001010111",
9613 => "001100110",
9614 => "001011011",
9615 => "001011101",
9616 => "001100101",
9617 => "001100110",
9618 => "001100000",
9619 => "001100100",
9620 => "001100011",
9621 => "001100111",
9622 => "001100110",
9623 => "001101010",
9624 => "001100111",
9625 => "001101011",
9626 => "001100010",
9627 => "001101000",
9628 => "001100111",
9629 => "001011100",
9630 => "001100011",
9631 => "001110011",
9632 => "001101010",
9633 => "001100111",
9634 => "001100010",
9635 => "001100001",
9636 => "001011111",
9637 => "001100010",
9638 => "001100011",
9639 => "001100010",
9640 => "001100111",
9641 => "001010110",
9642 => "001010111",
9643 => "001011100",
9644 => "001010101",
9645 => "001100010",
9646 => "001100000",
9647 => "001011001",
9648 => "001011100",
9649 => "001011110",
9650 => "001010010",
9651 => "001010010",
9652 => "001011001",
9653 => "001011001",
9654 => "001011011",
9655 => "001100101",
9656 => "001011101",
9657 => "001100000",
9658 => "001100001",
9659 => "001100001",
9660 => "001100000",
9661 => "001011010",
9662 => "001010101",
9663 => "001011000",
9664 => "001100001",
9665 => "001100010",
9666 => "001100100",
9667 => "001011101",
9668 => "001011011",
9669 => "001011000",
9670 => "001011100",
9671 => "001100000",
9672 => "001011111",
9673 => "001011101",
9674 => "001011010",
9675 => "001010110",
9676 => "001010110",
9677 => "001001011",
9678 => "000111110",
9679 => "001000001",
9680 => "001001101",
9681 => "001001011",
9682 => "001001100",
9683 => "001000110",
9684 => "001001011",
9685 => "001001001",
9686 => "001000101",
9687 => "001001011",
9688 => "001000110",
9689 => "000111010",
9690 => "001010000",
9691 => "001011010",
9692 => "001100000",
9693 => "001011110",
9694 => "001011010",
9695 => "001100010",
9696 => "001101100",
9697 => "001101000",
9698 => "001011110",
9699 => "001011111",
9700 => "001100110",
9701 => "001100100",
9702 => "001011011",
9703 => "001100011",
9704 => "001101111",
9705 => "001110101",
9706 => "001101011",
9707 => "001011000",
9708 => "001010011",
9709 => "001010110",
9710 => "001011000",
9711 => "001010001",
9712 => "001000111",
9713 => "001001011",
9714 => "001010001",
9715 => "001001100",
9716 => "001011010",
9717 => "001010100",
9718 => "001010100",
9719 => "001010000",
9720 => "001010001",
9721 => "001010011",
9722 => "001010011",
9723 => "001010111",
9724 => "001010101",
9725 => "001010100",
9726 => "001010111",
9727 => "001010011",
9728 => "001100100",
9729 => "001010110",
9730 => "001000110",
9731 => "001000101",
9732 => "001000001",
9733 => "001001100",
9734 => "001001000",
9735 => "001011110",
9736 => "001100101",
9737 => "001000011",
9738 => "001011000",
9739 => "001000101",
9740 => "001011001",
9741 => "001110011",
9742 => "001100110",
9743 => "001100100",
9744 => "001100110",
9745 => "001101101",
9746 => "001100100",
9747 => "001101000",
9748 => "001101001",
9749 => "001011111",
9750 => "001100100",
9751 => "001100101",
9752 => "001100100",
9753 => "001101010",
9754 => "001100101",
9755 => "001100101",
9756 => "001100111",
9757 => "001100111",
9758 => "001100101",
9759 => "001101101",
9760 => "001101011",
9761 => "001101110",
9762 => "001101000",
9763 => "001100111",
9764 => "001101100",
9765 => "001100101",
9766 => "001100100",
9767 => "001101110",
9768 => "001101101",
9769 => "001101100",
9770 => "001100101",
9771 => "001100101",
9772 => "001011101",
9773 => "001100000",
9774 => "001100000",
9775 => "001100010",
9776 => "001011111",
9777 => "001100000",
9778 => "001011010",
9779 => "001011101",
9780 => "001011000",
9781 => "001010110",
9782 => "001100111",
9783 => "001100101",
9784 => "001100011",
9785 => "001011011",
9786 => "001011001",
9787 => "001010110",
9788 => "001011110",
9789 => "001101000",
9790 => "001100100",
9791 => "001100000",
9792 => "001011110",
9793 => "001011100",
9794 => "001100000",
9795 => "001100100",
9796 => "001011101",
9797 => "001011100",
9798 => "001100010",
9799 => "001011101",
9800 => "001011111",
9801 => "001011101",
9802 => "001011100",
9803 => "001011001",
9804 => "001010111",
9805 => "001011001",
9806 => "001100011",
9807 => "001100010",
9808 => "001011100",
9809 => "001011001",
9810 => "001010111",
9811 => "001011001",
9812 => "001011001",
9813 => "001001011",
9814 => "001001110",
9815 => "001001000",
9816 => "001001001",
9817 => "000111100",
9818 => "001000001",
9819 => "001000100",
9820 => "001010101",
9821 => "001010110",
9822 => "001011110",
9823 => "001011100",
9824 => "001100001",
9825 => "001011111",
9826 => "001011001",
9827 => "001010011",
9828 => "001010011",
9829 => "001010001",
9830 => "001011000",
9831 => "001011000",
9832 => "001011101",
9833 => "001011001",
9834 => "001011010",
9835 => "001010100",
9836 => "001010001",
9837 => "001010001",
9838 => "001010110",
9839 => "001010110",
9840 => "001010010",
9841 => "001011001",
9842 => "001010111",
9843 => "001011001",
9844 => "001010101",
9845 => "001011001",
9846 => "001010110",
9847 => "001010010",
9848 => "001010111",
9849 => "001011011",
9850 => "001010100",
9851 => "001010110",
9852 => "001010110",
9853 => "001010100",
9854 => "001011001",
9855 => "001010100",
9856 => "001000110",
9857 => "000111110",
9858 => "001010001",
9859 => "000101111",
9860 => "001000101",
9861 => "001001000",
9862 => "001011000",
9863 => "000111010",
9864 => "000101010",
9865 => "000111101",
9866 => "000100101",
9867 => "000101011",
9868 => "001010100",
9869 => "001010111",
9870 => "001101011",
9871 => "001011111",
9872 => "001101000",
9873 => "001101010",
9874 => "001101101",
9875 => "001101010",
9876 => "001101001",
9877 => "001101000",
9878 => "001101110",
9879 => "001101110",
9880 => "001100101",
9881 => "001101110",
9882 => "001101101",
9883 => "001100111",
9884 => "001100010",
9885 => "001101001",
9886 => "001101000",
9887 => "001101011",
9888 => "001101101",
9889 => "001100000",
9890 => "001101001",
9891 => "001101010",
9892 => "001110001",
9893 => "001100101",
9894 => "001100011",
9895 => "001100100",
9896 => "001101000",
9897 => "001101011",
9898 => "001100110",
9899 => "001100110",
9900 => "001100110",
9901 => "001100011",
9902 => "001011111",
9903 => "001100111",
9904 => "001100101",
9905 => "001101010",
9906 => "001100001",
9907 => "001011111",
9908 => "001100000",
9909 => "001100010",
9910 => "001011111",
9911 => "001010110",
9912 => "001011110",
9913 => "001011101",
9914 => "001100000",
9915 => "001011110",
9916 => "001011110",
9917 => "001011000",
9918 => "001001111",
9919 => "001110101",
9920 => "001101101",
9921 => "001100111",
9922 => "001100111",
9923 => "001100101",
9924 => "001011101",
9925 => "001011100",
9926 => "001101001",
9927 => "001100110",
9928 => "001100001",
9929 => "001011100",
9930 => "001011100",
9931 => "001100011",
9932 => "001100010",
9933 => "001100101",
9934 => "001011111",
9935 => "001010111",
9936 => "001011001",
9937 => "001010110",
9938 => "001011011",
9939 => "001010011",
9940 => "001010111",
9941 => "001010110",
9942 => "001010000",
9943 => "001011000",
9944 => "001010001",
9945 => "001100101",
9946 => "001011000",
9947 => "001000010",
9948 => "001000010",
9949 => "001000111",
9950 => "001001111",
9951 => "001010100",
9952 => "001010101",
9953 => "001010100",
9954 => "001010111",
9955 => "001001111",
9956 => "001010010",
9957 => "001010011",
9958 => "001011001",
9959 => "001011011",
9960 => "001011101",
9961 => "001010111",
9962 => "001010110",
9963 => "001010111",
9964 => "001010110",
9965 => "001011011",
9966 => "001011011",
9967 => "001010100",
9968 => "001010011",
9969 => "001010010",
9970 => "001010100",
9971 => "001010011",
9972 => "001010001",
9973 => "001010110",
9974 => "001010000",
9975 => "001010110",
9976 => "001010110",
9977 => "001010010",
9978 => "001011010",
9979 => "001011001",
9980 => "001010100",
9981 => "001010010",
9982 => "001011000",
9983 => "001010110",
9984 => "000110001",
9985 => "000101001",
9986 => "001001011",
9987 => "001010011",
9988 => "001001011",
9989 => "001001010",
9990 => "001010101",
9991 => "001010100",
9992 => "000111001",
9993 => "001010110",
9994 => "000101111",
9995 => "001001100",
9996 => "001000111",
9997 => "001010111",
9998 => "001110000",
9999 => "001100011",
10000 => "001100000",
10001 => "001100101",
10002 => "001100001",
10003 => "001100100",
10004 => "001100110",
10005 => "001100101",
10006 => "001101011",
10007 => "001101011",
10008 => "001101000",
10009 => "001101000",
10010 => "001110001",
10011 => "001110001",
10012 => "001110010",
10013 => "001110000",
10014 => "001110010",
10015 => "001101101",
10016 => "001110011",
10017 => "001110100",
10018 => "001101010",
10019 => "001101011",
10020 => "001101101",
10021 => "001110000",
10022 => "001100110",
10023 => "001100111",
10024 => "001100100",
10025 => "001101100",
10026 => "001101001",
10027 => "001101001",
10028 => "001100101",
10029 => "001101111",
10030 => "001101011",
10031 => "001101000",
10032 => "001100110",
10033 => "001101001",
10034 => "001100110",
10035 => "001101010",
10036 => "001100100",
10037 => "001100111",
10038 => "001100001",
10039 => "001011010",
10040 => "001010001",
10041 => "001001101",
10042 => "001010100",
10043 => "001100001",
10044 => "001100001",
10045 => "001101001",
10046 => "001100110",
10047 => "001011000",
10048 => "001011100",
10049 => "001100100",
10050 => "001100110",
10051 => "001100110",
10052 => "001010110",
10053 => "001011101",
10054 => "001100001",
10055 => "001100100",
10056 => "001100110",
10057 => "001011111",
10058 => "001011101",
10059 => "001011011",
10060 => "001011011",
10061 => "001100011",
10062 => "001100000",
10063 => "001100010",
10064 => "001100011",
10065 => "001100001",
10066 => "001011010",
10067 => "001011010",
10068 => "001011000",
10069 => "001001111",
10070 => "001010100",
10071 => "001010100",
10072 => "001011001",
10073 => "001010010",
10074 => "001010100",
10075 => "001010110",
10076 => "001010100",
10077 => "001010001",
10078 => "001011001",
10079 => "001011010",
10080 => "001010101",
10081 => "001011010",
10082 => "001011000",
10083 => "001010101",
10084 => "001010101",
10085 => "001010110",
10086 => "001011010",
10087 => "001011001",
10088 => "001011000",
10089 => "001010100",
10090 => "001011001",
10091 => "001010110",
10092 => "001010011",
10093 => "001010001",
10094 => "001010010",
10095 => "001010101",
10096 => "001010110",
10097 => "001010111",
10098 => "001010100",
10099 => "001010110",
10100 => "001011010",
10101 => "001010111",
10102 => "001010111",
10103 => "001011001",
10104 => "001010111",
10105 => "001010110",
10106 => "001010100",
10107 => "001011000",
10108 => "001010101",
10109 => "001011000",
10110 => "001011000",
10111 => "001011010",
10112 => "001011011",
10113 => "000110001",
10114 => "000111111",
10115 => "000111011",
10116 => "001000010",
10117 => "001001101",
10118 => "001000110",
10119 => "000111000",
10120 => "000111100",
10121 => "001000101",
10122 => "001001100",
10123 => "001010010",
10124 => "001011000",
10125 => "001010000",
10126 => "001101101",
10127 => "001100010",
10128 => "001100000",
10129 => "001011110",
10130 => "001101101",
10131 => "001101010",
10132 => "001100110",
10133 => "001100110",
10134 => "001011010",
10135 => "001100001",
10136 => "001100010",
10137 => "001100100",
10138 => "001100110",
10139 => "001100001",
10140 => "001100111",
10141 => "001101010",
10142 => "001100111",
10143 => "001101001",
10144 => "001101000",
10145 => "001100000",
10146 => "001011100",
10147 => "001101011",
10148 => "001101000",
10149 => "001100110",
10150 => "001100111",
10151 => "001100111",
10152 => "001101110",
10153 => "001101000",
10154 => "001100111",
10155 => "001101010",
10156 => "001110000",
10157 => "001101101",
10158 => "001110001",
10159 => "001101110",
10160 => "001101011",
10161 => "001100101",
10162 => "001100011",
10163 => "001101101",
10164 => "001100111",
10165 => "001101000",
10166 => "001100110",
10167 => "001100010",
10168 => "001011111",
10169 => "001100000",
10170 => "001011010",
10171 => "001010111",
10172 => "001011100",
10173 => "001011010",
10174 => "001100000",
10175 => "001011010",
10176 => "001011000",
10177 => "001011100",
10178 => "001101000",
10179 => "001101100",
10180 => "001011100",
10181 => "001011000",
10182 => "001100011",
10183 => "001100011",
10184 => "001100001",
10185 => "001011011",
10186 => "001100110",
10187 => "001011111",
10188 => "001011100",
10189 => "001011000",
10190 => "001011011",
10191 => "001011101",
10192 => "001011001",
10193 => "001011100",
10194 => "001011101",
10195 => "001011110",
10196 => "001100001",
10197 => "001100001",
10198 => "001011100",
10199 => "001011010",
10200 => "001010010",
10201 => "001011100",
10202 => "001100011",
10203 => "001011011",
10204 => "001011110",
10205 => "001011000",
10206 => "001010110",
10207 => "001011010",
10208 => "001011101",
10209 => "001100011",
10210 => "001110110",
10211 => "001011110",
10212 => "001011001",
10213 => "001011011",
10214 => "001011011",
10215 => "001011110",
10216 => "001011101",
10217 => "001011010",
10218 => "001011011",
10219 => "001011010",
10220 => "001011001",
10221 => "001011100",
10222 => "001011001",
10223 => "001011101",
10224 => "001011100",
10225 => "001010101",
10226 => "001010100",
10227 => "001010000",
10228 => "001010011",
10229 => "001011001",
10230 => "001010101",
10231 => "001010100",
10232 => "001010100",
10233 => "001010101",
10234 => "001010010",
10235 => "001001110",
10236 => "001010100",
10237 => "001010111",
10238 => "001010001",
10239 => "001010101",
10240 => "001010001",
10241 => "001001110",
10242 => "000111000",
10243 => "000110101",
10244 => "001001101",
10245 => "001001100",
10246 => "001000110",
10247 => "001001011",
10248 => "000101011",
10249 => "000110011",
10250 => "001001010",
10251 => "001011001",
10252 => "001101000",
10253 => "001011111",
10254 => "001101001",
10255 => "001011010",
10256 => "001011001",
10257 => "001100101",
10258 => "001100111",
10259 => "001101010",
10260 => "001101011",
10261 => "001101110",
10262 => "001101101",
10263 => "001100111",
10264 => "001101000",
10265 => "001101000",
10266 => "001100110",
10267 => "001100111",
10268 => "001011111",
10269 => "001011111",
10270 => "001100010",
10271 => "001100010",
10272 => "001101001",
10273 => "001101001",
10274 => "001100101",
10275 => "001101010",
10276 => "001101001",
10277 => "001100100",
10278 => "001101001",
10279 => "001101111",
10280 => "001110000",
10281 => "001101100",
10282 => "001101101",
10283 => "001110001",
10284 => "001101100",
10285 => "001101011",
10286 => "001101010",
10287 => "001100110",
10288 => "001100111",
10289 => "001101110",
10290 => "001101101",
10291 => "001101011",
10292 => "001101000",
10293 => "001101001",
10294 => "001100101",
10295 => "001101001",
10296 => "001100100",
10297 => "001011111",
10298 => "001100100",
10299 => "001100001",
10300 => "001100010",
10301 => "001011110",
10302 => "001100100",
10303 => "001100001",
10304 => "001100100",
10305 => "001011111",
10306 => "001100111",
10307 => "001101000",
10308 => "001101000",
10309 => "001101000",
10310 => "001101101",
10311 => "001100110",
10312 => "001100111",
10313 => "001100110",
10314 => "001100010",
10315 => "001100100",
10316 => "001011100",
10317 => "001011011",
10318 => "001011110",
10319 => "001011111",
10320 => "001011111",
10321 => "001011011",
10322 => "001100000",
10323 => "001100101",
10324 => "001100101",
10325 => "001100111",
10326 => "001100100",
10327 => "001100100",
10328 => "001100011",
10329 => "001011111",
10330 => "001011001",
10331 => "001010000",
10332 => "001010110",
10333 => "001011111",
10334 => "001100101",
10335 => "001100001",
10336 => "001100010",
10337 => "001100011",
10338 => "001011111",
10339 => "001100001",
10340 => "001011101",
10341 => "001011111",
10342 => "001011010",
10343 => "001011010",
10344 => "001010101",
10345 => "001011101",
10346 => "001011101",
10347 => "001011010",
10348 => "001010100",
10349 => "001010010",
10350 => "001010010",
10351 => "001010011",
10352 => "001010110",
10353 => "001010111",
10354 => "001010101",
10355 => "001011001",
10356 => "001011001",
10357 => "001011010",
10358 => "001011000",
10359 => "001010100",
10360 => "001010110",
10361 => "001010111",
10362 => "001011010",
10363 => "001011101",
10364 => "001011100",
10365 => "001010110",
10366 => "001010100",
10367 => "001010101",
10368 => "001000100",
10369 => "001010001",
10370 => "000111000",
10371 => "000111010",
10372 => "000101101",
10373 => "001001010",
10374 => "001000001",
10375 => "001001101",
10376 => "001010000",
10377 => "000111011",
10378 => "001001111",
10379 => "001010000",
10380 => "001011100",
10381 => "001010001",
10382 => "001100010",
10383 => "001100010",
10384 => "001100000",
10385 => "001011101",
10386 => "001100010",
10387 => "001011111",
10388 => "001011011",
10389 => "001100110",
10390 => "001011100",
10391 => "001011000",
10392 => "001100001",
10393 => "001011101",
10394 => "001101011",
10395 => "001101001",
10396 => "001101001",
10397 => "001101100",
10398 => "001101001",
10399 => "001100111",
10400 => "001101110",
10401 => "001100111",
10402 => "001100111",
10403 => "001011001",
10404 => "001101101",
10405 => "001100111",
10406 => "001011110",
10407 => "001010101",
10408 => "001100001",
10409 => "001101110",
10410 => "001101100",
10411 => "001101010",
10412 => "001100111",
10413 => "001101011",
10414 => "001101000",
10415 => "001101001",
10416 => "001101000",
10417 => "001101010",
10418 => "001110111",
10419 => "001101110",
10420 => "001101010",
10421 => "001101110",
10422 => "001101100",
10423 => "001101110",
10424 => "001101011",
10425 => "001101001",
10426 => "001110100",
10427 => "001101111",
10428 => "001110000",
10429 => "001100111",
10430 => "001100110",
10431 => "001100110",
10432 => "001100110",
10433 => "001101001",
10434 => "001101010",
10435 => "001101101",
10436 => "001100101",
10437 => "001101000",
10438 => "001101111",
10439 => "001101001",
10440 => "001101010",
10441 => "001101010",
10442 => "001101000",
10443 => "001100000",
10444 => "001011111",
10445 => "001100011",
10446 => "001101000",
10447 => "001100101",
10448 => "001100011",
10449 => "001100100",
10450 => "001100110",
10451 => "001100111",
10452 => "001100000",
10453 => "001100011",
10454 => "001011111",
10455 => "001011010",
10456 => "001100011",
10457 => "001010011",
10458 => "001010101",
10459 => "001001110",
10460 => "001001111",
10461 => "001011011",
10462 => "001011101",
10463 => "001011101",
10464 => "001011010",
10465 => "001011011",
10466 => "001011101",
10467 => "001010111",
10468 => "001011001",
10469 => "001011100",
10470 => "001100010",
10471 => "001011100",
10472 => "001011111",
10473 => "001011110",
10474 => "001011100",
10475 => "001010011",
10476 => "001011001",
10477 => "001011101",
10478 => "001100000",
10479 => "001100001",
10480 => "001011110",
10481 => "001011001",
10482 => "001011100",
10483 => "001011011",
10484 => "001011111",
10485 => "001011100",
10486 => "001011011",
10487 => "001011110",
10488 => "001011000",
10489 => "001001101",
10490 => "001001110",
10491 => "001010110",
10492 => "001010011",
10493 => "001010001",
10494 => "001011101",
10495 => "001011001",
10496 => "000111001",
10497 => "001010011",
10498 => "000101111",
10499 => "000101011",
10500 => "000100111",
10501 => "000111101",
10502 => "001000110",
10503 => "001001011",
10504 => "001011110",
10505 => "001010011",
10506 => "001010010",
10507 => "001001011",
10508 => "001100110",
10509 => "001100101",
10510 => "001100011",
10511 => "001101001",
10512 => "001100001",
10513 => "001011100",
10514 => "001100101",
10515 => "001011000",
10516 => "001100101",
10517 => "001011111",
10518 => "001011001",
10519 => "001011011",
10520 => "001011110",
10521 => "001101000",
10522 => "001011000",
10523 => "001011111",
10524 => "001100110",
10525 => "001100010",
10526 => "001101010",
10527 => "001101110",
10528 => "001101111",
10529 => "001101010",
10530 => "001101011",
10531 => "001101001",
10532 => "001101110",
10533 => "001101101",
10534 => "001101011",
10535 => "001100011",
10536 => "001100010",
10537 => "001100011",
10538 => "001011111",
10539 => "001101001",
10540 => "001011111",
10541 => "001100110",
10542 => "001100111",
10543 => "001101011",
10544 => "001101000",
10545 => "001100110",
10546 => "001110011",
10547 => "001110111",
10548 => "001110000",
10549 => "001110001",
10550 => "001110101",
10551 => "001101001",
10552 => "001100111",
10553 => "001110001",
10554 => "001111001",
10555 => "001110101",
10556 => "001100110",
10557 => "001101101",
10558 => "001100101",
10559 => "001101000",
10560 => "001100010",
10561 => "001101110",
10562 => "001101010",
10563 => "001110001",
10564 => "001110010",
10565 => "001110010",
10566 => "001101110",
10567 => "001111101",
10568 => "001110000",
10569 => "001101110",
10570 => "001110000",
10571 => "001101110",
10572 => "001110010",
10573 => "001110000",
10574 => "001100100",
10575 => "001101010",
10576 => "001101001",
10577 => "001100110",
10578 => "001011111",
10579 => "001011001",
10580 => "001010111",
10581 => "001100101",
10582 => "001100010",
10583 => "001100100",
10584 => "001011101",
10585 => "001011111",
10586 => "001011100",
10587 => "001011000",
10588 => "001100011",
10589 => "001100001",
10590 => "001011101",
10591 => "001100101",
10592 => "001100110",
10593 => "001100000",
10594 => "001100000",
10595 => "001011001",
10596 => "001011100",
10597 => "001011111",
10598 => "001011101",
10599 => "001011101",
10600 => "001011001",
10601 => "001001110",
10602 => "001011100",
10603 => "001100000",
10604 => "001100010",
10605 => "001100000",
10606 => "001100011",
10607 => "001011111",
10608 => "001011111",
10609 => "001100001",
10610 => "001011100",
10611 => "001011100",
10612 => "001011010",
10613 => "001010011",
10614 => "001010100",
10615 => "001010100",
10616 => "001011001",
10617 => "001011000",
10618 => "001010100",
10619 => "001011110",
10620 => "001010001",
10621 => "001011001",
10622 => "001011000",
10623 => "001011000",
10624 => "001010001",
10625 => "001010110",
10626 => "000111110",
10627 => "000011100",
10628 => "000101000",
10629 => "001000000",
10630 => "000101101",
10631 => "001001011",
10632 => "001100010",
10633 => "000110100",
10634 => "001001010",
10635 => "001011100",
10636 => "001100011",
10637 => "001011011",
10638 => "001010110",
10639 => "001011011",
10640 => "001100101",
10641 => "001100010",
10642 => "001011011",
10643 => "001001010",
10644 => "001100101",
10645 => "001101001",
10646 => "001011010",
10647 => "001100011",
10648 => "001010111",
10649 => "001101101",
10650 => "001101101",
10651 => "001011101",
10652 => "001100010",
10653 => "001100110",
10654 => "001011001",
10655 => "001011001",
10656 => "001100011",
10657 => "001100010",
10658 => "001100011",
10659 => "001101101",
10660 => "001100101",
10661 => "001101000",
10662 => "001110001",
10663 => "001101000",
10664 => "001101001",
10665 => "001100000",
10666 => "001100110",
10667 => "001101001",
10668 => "001101000",
10669 => "001101000",
10670 => "001101001",
10671 => "001101101",
10672 => "001110011",
10673 => "001101011",
10674 => "001101001",
10675 => "001100111",
10676 => "001101101",
10677 => "001100111",
10678 => "001100111",
10679 => "001101000",
10680 => "001101100",
10681 => "001110010",
10682 => "001111000",
10683 => "001110001",
10684 => "001110010",
10685 => "001101010",
10686 => "001101010",
10687 => "001010111",
10688 => "001010010",
10689 => "001100101",
10690 => "001100101",
10691 => "001011111",
10692 => "001101110",
10693 => "001101110",
10694 => "001100100",
10695 => "001101000",
10696 => "001101110",
10697 => "001110111",
10698 => "001110111",
10699 => "001110101",
10700 => "001110011",
10701 => "001111010",
10702 => "001111001",
10703 => "001110011",
10704 => "001110110",
10705 => "001110001",
10706 => "001110010",
10707 => "001101000",
10708 => "001101100",
10709 => "001110111",
10710 => "001101101",
10711 => "001101111",
10712 => "001101110",
10713 => "001100011",
10714 => "001011011",
10715 => "001100111",
10716 => "001101101",
10717 => "001101010",
10718 => "001101000",
10719 => "001100101",
10720 => "001011101",
10721 => "001011010",
10722 => "001010101",
10723 => "001010100",
10724 => "001011111",
10725 => "001100110",
10726 => "001100000",
10727 => "001100100",
10728 => "001100001",
10729 => "001011110",
10730 => "001010101",
10731 => "001011101",
10732 => "001011000",
10733 => "001011110",
10734 => "001011111",
10735 => "001011100",
10736 => "001011010",
10737 => "001011000",
10738 => "001100010",
10739 => "001100010",
10740 => "001011111",
10741 => "001011011",
10742 => "001100010",
10743 => "001101110",
10744 => "001101000",
10745 => "001011100",
10746 => "001101001",
10747 => "001100001",
10748 => "001100011",
10749 => "001010011",
10750 => "001001101",
10751 => "001010111",
10752 => "000100110",
10753 => "000111011",
10754 => "000110000",
10755 => "000110011",
10756 => "000101100",
10757 => "001001000",
10758 => "001010111",
10759 => "000111011",
10760 => "001011111",
10761 => "001100111",
10762 => "001001101",
10763 => "001001001",
10764 => "001100010",
10765 => "001100110",
10766 => "001100100",
10767 => "001100101",
10768 => "001100101",
10769 => "001011110",
10770 => "001010101",
10771 => "001101101",
10772 => "001011100",
10773 => "001010000",
10774 => "001010110",
10775 => "001010000",
10776 => "001100101",
10777 => "001011110",
10778 => "001011101",
10779 => "001011011",
10780 => "001011010",
10781 => "001011100",
10782 => "001010110",
10783 => "001010100",
10784 => "001010110",
10785 => "001100001",
10786 => "001100101",
10787 => "001010110",
10788 => "001010101",
10789 => "001011011",
10790 => "001010010",
10791 => "001101100",
10792 => "001100010",
10793 => "001010011",
10794 => "001010010",
10795 => "001011010",
10796 => "001100001",
10797 => "001100111",
10798 => "001101000",
10799 => "001100000",
10800 => "001011111",
10801 => "001100100",
10802 => "001101111",
10803 => "001101001",
10804 => "001100110",
10805 => "001101111",
10806 => "001100100",
10807 => "001101001",
10808 => "001100111",
10809 => "001011010",
10810 => "001101010",
10811 => "001101101",
10812 => "001101101",
10813 => "001110001",
10814 => "001101101",
10815 => "001101011",
10816 => "001101100",
10817 => "001100101",
10818 => "001101100",
10819 => "001101011",
10820 => "001100101",
10821 => "001101101",
10822 => "001100101",
10823 => "001100111",
10824 => "001101111",
10825 => "001100101",
10826 => "001101101",
10827 => "001101111",
10828 => "001110010",
10829 => "001110110",
10830 => "001110011",
10831 => "001110101",
10832 => "001110011",
10833 => "001110001",
10834 => "001110010",
10835 => "001110000",
10836 => "001110000",
10837 => "001110101",
10838 => "001101111",
10839 => "001100100",
10840 => "001101011",
10841 => "001100110",
10842 => "001100010",
10843 => "001101010",
10844 => "001011101",
10845 => "001100111",
10846 => "001100001",
10847 => "001101101",
10848 => "001110000",
10849 => "001100001",
10850 => "001100000",
10851 => "001011001",
10852 => "001011011",
10853 => "001100001",
10854 => "001011001",
10855 => "001010011",
10856 => "001011110",
10857 => "001100111",
10858 => "001100001",
10859 => "001100100",
10860 => "001011100",
10861 => "001010110",
10862 => "001011010",
10863 => "001011101",
10864 => "001011001",
10865 => "001011010",
10866 => "001010000",
10867 => "001001001",
10868 => "001001110",
10869 => "001001110",
10870 => "001011101",
10871 => "001011000",
10872 => "001100001",
10873 => "001010011",
10874 => "001001010",
10875 => "001001001",
10876 => "001011100",
10877 => "001100000",
10878 => "001100011",
10879 => "001011011",
10880 => "000100100",
10881 => "000011101",
10882 => "000100001",
10883 => "000111100",
10884 => "000011111",
10885 => "000011111",
10886 => "001011011",
10887 => "001011011",
10888 => "001011011",
10889 => "001101110",
10890 => "001011110",
10891 => "001010001",
10892 => "001011110",
10893 => "001100111",
10894 => "001011001",
10895 => "001010000",
10896 => "001011101",
10897 => "001011001",
10898 => "001101000",
10899 => "001101101",
10900 => "001100001",
10901 => "001100010",
10902 => "001100001",
10903 => "001011110",
10904 => "001011011",
10905 => "001010000",
10906 => "001011001",
10907 => "001100100",
10908 => "001101011",
10909 => "001100110",
10910 => "001100001",
10911 => "001100000",
10912 => "001100000",
10913 => "001100111",
10914 => "001011101",
10915 => "001011100",
10916 => "001011111",
10917 => "001100010",
10918 => "001011011",
10919 => "001011111",
10920 => "001100100",
10921 => "001101010",
10922 => "001100100",
10923 => "001100101",
10924 => "001100010",
10925 => "001011111",
10926 => "001100001",
10927 => "001100011",
10928 => "001101000",
10929 => "001100100",
10930 => "001101110",
10931 => "001101001",
10932 => "001100110",
10933 => "001101001",
10934 => "001100111",
10935 => "001011111",
10936 => "001101000",
10937 => "001100101",
10938 => "001011110",
10939 => "001001111",
10940 => "001100000",
10941 => "001110010",
10942 => "001110001",
10943 => "001100110",
10944 => "001100111",
10945 => "001101101",
10946 => "001100101",
10947 => "001100111",
10948 => "001011110",
10949 => "001101001",
10950 => "001110101",
10951 => "001110010",
10952 => "001101111",
10953 => "001100110",
10954 => "001110001",
10955 => "001101010",
10956 => "001101011",
10957 => "001101011",
10958 => "001110001",
10959 => "001110111",
10960 => "001111010",
10961 => "001110001",
10962 => "001110101",
10963 => "001110010",
10964 => "001111001",
10965 => "001101101",
10966 => "001101110",
10967 => "001110000",
10968 => "001101000",
10969 => "001100001",
10970 => "001101010",
10971 => "001100101",
10972 => "001100010",
10973 => "001011101",
10974 => "001100101",
10975 => "001101000",
10976 => "001100000",
10977 => "001100100",
10978 => "001100000",
10979 => "001011011",
10980 => "001011101",
10981 => "001001110",
10982 => "001011110",
10983 => "001011011",
10984 => "001010110",
10985 => "001011101",
10986 => "001100010",
10987 => "001100101",
10988 => "001100010",
10989 => "001011101",
10990 => "001011000",
10991 => "001100100",
10992 => "001011011",
10993 => "001010100",
10994 => "001010111",
10995 => "001011000",
10996 => "001011101",
10997 => "001011001",
10998 => "001010001",
10999 => "001010100",
11000 => "001011010",
11001 => "001011000",
11002 => "001010100",
11003 => "001011110",
11004 => "001100010",
11005 => "001100000",
11006 => "001100001",
11007 => "001011100",
11008 => "000011100",
11009 => "000010111",
11010 => "000010110",
11011 => "000011011",
11012 => "000100000",
11013 => "000111001",
11014 => "000110011",
11015 => "000110100",
11016 => "001011111",
11017 => "001011011",
11018 => "001000100",
11019 => "001000001",
11020 => "001101111",
11021 => "001101001",
11022 => "001010111",
11023 => "001100010",
11024 => "001101101",
11025 => "001101000",
11026 => "001101110",
11027 => "001100011",
11028 => "001011010",
11029 => "001100111",
11030 => "001011111",
11031 => "001101100",
11032 => "001100101",
11033 => "001101000",
11034 => "001101111",
11035 => "001101111",
11036 => "001101110",
11037 => "001100110",
11038 => "001101011",
11039 => "001101000",
11040 => "001100100",
11041 => "001100111",
11042 => "001101111",
11043 => "001100111",
11044 => "001100000",
11045 => "001011101",
11046 => "001011010",
11047 => "001100101",
11048 => "001100100",
11049 => "001100101",
11050 => "001100000",
11051 => "001101001",
11052 => "001101000",
11053 => "001101110",
11054 => "001101000",
11055 => "001101010",
11056 => "001101011",
11057 => "001100101",
11058 => "001100100",
11059 => "001011111",
11060 => "001100010",
11061 => "001011010",
11062 => "001010111",
11063 => "001100100",
11064 => "001100011",
11065 => "001101101",
11066 => "001100100",
11067 => "001100100",
11068 => "001100010",
11069 => "001101000",
11070 => "001101100",
11071 => "001101011",
11072 => "001101011",
11073 => "001101110",
11074 => "001110011",
11075 => "001101100",
11076 => "001100101",
11077 => "001011111",
11078 => "001110000",
11079 => "001101001",
11080 => "001101110",
11081 => "001101110",
11082 => "001110001",
11083 => "001101010",
11084 => "001101001",
11085 => "001110100",
11086 => "001110000",
11087 => "001110101",
11088 => "001100001",
11089 => "001100100",
11090 => "001101010",
11091 => "001101000",
11092 => "001110010",
11093 => "001101110",
11094 => "001110001",
11095 => "001110000",
11096 => "001110000",
11097 => "001101011",
11098 => "001101011",
11099 => "001110010",
11100 => "001101100",
11101 => "001101000",
11102 => "001011000",
11103 => "001100100",
11104 => "001110000",
11105 => "001100111",
11106 => "001011100",
11107 => "001010001",
11108 => "001010101",
11109 => "001010011",
11110 => "001011000",
11111 => "001010111",
11112 => "001001110",
11113 => "001001100",
11114 => "001001110",
11115 => "001011011",
11116 => "001010011",
11117 => "001010101",
11118 => "001010011",
11119 => "001010001",
11120 => "001010110",
11121 => "001011010",
11122 => "001011011",
11123 => "001011001",
11124 => "001011101",
11125 => "001010111",
11126 => "001100000",
11127 => "001011100",
11128 => "001011100",
11129 => "001010111",
11130 => "001001110",
11131 => "001010101",
11132 => "001010011",
11133 => "001010101",
11134 => "001011010",
11135 => "001011111",
11136 => "001010001",
11137 => "001011001",
11138 => "001110111",
11139 => "000101101",
11140 => "001000001",
11141 => "001000000",
11142 => "000101011",
11143 => "001000000",
11144 => "001010001",
11145 => "001010001",
11146 => "001010100",
11147 => "001101010",
11148 => "001011010",
11149 => "001011000",
11150 => "001100011",
11151 => "001010100",
11152 => "001101010",
11153 => "001011001",
11154 => "001101000",
11155 => "001100100",
11156 => "001110001",
11157 => "001110001",
11158 => "001100011",
11159 => "001100001",
11160 => "001011010",
11161 => "001011111",
11162 => "001100011",
11163 => "001100010",
11164 => "001100111",
11165 => "001110001",
11166 => "001101000",
11167 => "001100101",
11168 => "001101101",
11169 => "001101011",
11170 => "001101101",
11171 => "001101010",
11172 => "001101000",
11173 => "001100101",
11174 => "001100001",
11175 => "001100101",
11176 => "001011101",
11177 => "001100011",
11178 => "001100101",
11179 => "001011011",
11180 => "001011100",
11181 => "001011011",
11182 => "001010110",
11183 => "001101010",
11184 => "001100011",
11185 => "001100101",
11186 => "001011111",
11187 => "001011011",
11188 => "001011000",
11189 => "001100010",
11190 => "001100100",
11191 => "001011111",
11192 => "001011111",
11193 => "001100110",
11194 => "001010101",
11195 => "001011111",
11196 => "001100111",
11197 => "001100111",
11198 => "001101101",
11199 => "001101001",
11200 => "001100100",
11201 => "001101110",
11202 => "001100011",
11203 => "001011111",
11204 => "001101110",
11205 => "001110000",
11206 => "001101000",
11207 => "001110010",
11208 => "001101010",
11209 => "001100111",
11210 => "001101101",
11211 => "001101111",
11212 => "001100111",
11213 => "001110001",
11214 => "001101011",
11215 => "001101101",
11216 => "001110000",
11217 => "001100100",
11218 => "001111010",
11219 => "001101100",
11220 => "001110100",
11221 => "001110000",
11222 => "001110111",
11223 => "001101111",
11224 => "001110010",
11225 => "001101100",
11226 => "001101100",
11227 => "001101010",
11228 => "001111001",
11229 => "001100011",
11230 => "001101010",
11231 => "001100100",
11232 => "001101101",
11233 => "001101010",
11234 => "001100101",
11235 => "001100110",
11236 => "001100110",
11237 => "001011111",
11238 => "001101000",
11239 => "001011100",
11240 => "001011011",
11241 => "001010111",
11242 => "001011000",
11243 => "001100001",
11244 => "001011110",
11245 => "001010111",
11246 => "001011001",
11247 => "001011110",
11248 => "001011000",
11249 => "001010010",
11250 => "001010010",
11251 => "001100011",
11252 => "001011010",
11253 => "001011001",
11254 => "001010000",
11255 => "001010111",
11256 => "001010011",
11257 => "001100001",
11258 => "001011000",
11259 => "001011111",
11260 => "001011111",
11261 => "001011100",
11262 => "001100001",
11263 => "001010011",
11264 => "001001100",
11265 => "001001000",
11266 => "000110000",
11267 => "000111101",
11268 => "001000001",
11269 => "000111100",
11270 => "001100100",
11271 => "001000010",
11272 => "000111000",
11273 => "001010101",
11274 => "001100111",
11275 => "001001110",
11276 => "001000100",
11277 => "001000001",
11278 => "001110101",
11279 => "001010110",
11280 => "001011101",
11281 => "001111011",
11282 => "001100111",
11283 => "001101100",
11284 => "001100111",
11285 => "001110000",
11286 => "001100101",
11287 => "001100110",
11288 => "001100011",
11289 => "001011100",
11290 => "001100111",
11291 => "001100100",
11292 => "001101000",
11293 => "001011110",
11294 => "001011011",
11295 => "001100010",
11296 => "001100101",
11297 => "001011111",
11298 => "001101001",
11299 => "001101011",
11300 => "001101100",
11301 => "001101001",
11302 => "001101010",
11303 => "001100111",
11304 => "001100001",
11305 => "001100000",
11306 => "001101010",
11307 => "001101101",
11308 => "001100011",
11309 => "001011010",
11310 => "001010011",
11311 => "001010010",
11312 => "001010111",
11313 => "001100010",
11314 => "001011011",
11315 => "001100001",
11316 => "001010110",
11317 => "001011000",
11318 => "001101010",
11319 => "001100101",
11320 => "001100110",
11321 => "001100101",
11322 => "001100000",
11323 => "001100010",
11324 => "001100100",
11325 => "001110000",
11326 => "001100110",
11327 => "001101011",
11328 => "001101111",
11329 => "001101110",
11330 => "001110000",
11331 => "001110001",
11332 => "001101010",
11333 => "001101100",
11334 => "001110001",
11335 => "001101010",
11336 => "001101011",
11337 => "001101010",
11338 => "001101001",
11339 => "001110000",
11340 => "001101111",
11341 => "001110000",
11342 => "001101110",
11343 => "001101111",
11344 => "001101100",
11345 => "001100110",
11346 => "001101101",
11347 => "001101100",
11348 => "001110010",
11349 => "001101011",
11350 => "001101010",
11351 => "001101100",
11352 => "001110101",
11353 => "001101101",
11354 => "001110001",
11355 => "001100110",
11356 => "001110011",
11357 => "001101101",
11358 => "001101001",
11359 => "001100110",
11360 => "001101000",
11361 => "001110000",
11362 => "001101111",
11363 => "001101011",
11364 => "001101101",
11365 => "001100010",
11366 => "001100110",
11367 => "001100000",
11368 => "001100100",
11369 => "001011010",
11370 => "001010110",
11371 => "001011000",
11372 => "001100011",
11373 => "001100000",
11374 => "001010010",
11375 => "001010011",
11376 => "001100010",
11377 => "001011001",
11378 => "001011000",
11379 => "001010001",
11380 => "001001110",
11381 => "001011101",
11382 => "001010100",
11383 => "001011101",
11384 => "001010101",
11385 => "001011011",
11386 => "001010111",
11387 => "001011000",
11388 => "001011001",
11389 => "001100000",
11390 => "001011001",
11391 => "001011110",
11392 => "001010001",
11393 => "001001110",
11394 => "000010111",
11395 => "000101110",
11396 => "001000100",
11397 => "001000010",
11398 => "001000011",
11399 => "001001010",
11400 => "001011101",
11401 => "000111010",
11402 => "001000001",
11403 => "001001100",
11404 => "001000001",
11405 => "001000010",
11406 => "001011010",
11407 => "001001001",
11408 => "000111001",
11409 => "001011100",
11410 => "001110010",
11411 => "001101100",
11412 => "001101000",
11413 => "001101001",
11414 => "001100110",
11415 => "001010110",
11416 => "001001010",
11417 => "001001110",
11418 => "001000110",
11419 => "001001111",
11420 => "001100010",
11421 => "001100000",
11422 => "001100011",
11423 => "001101110",
11424 => "001100010",
11425 => "001100100",
11426 => "001100101",
11427 => "001011101",
11428 => "001011111",
11429 => "001100011",
11430 => "001101001",
11431 => "001100110",
11432 => "001101000",
11433 => "001100001",
11434 => "001100001",
11435 => "001100101",
11436 => "001100111",
11437 => "001101011",
11438 => "001100110",
11439 => "001100000",
11440 => "001100110",
11441 => "001101000",
11442 => "001100010",
11443 => "001011101",
11444 => "001100001",
11445 => "001100001",
11446 => "001010001",
11447 => "001010001",
11448 => "001010010",
11449 => "001101101",
11450 => "001100001",
11451 => "001100000",
11452 => "001011110",
11453 => "001100110",
11454 => "001101101",
11455 => "001101100",
11456 => "001101100",
11457 => "001101001",
11458 => "001101111",
11459 => "001100111",
11460 => "001101011",
11461 => "001101101",
11462 => "001101000",
11463 => "001101100",
11464 => "001110000",
11465 => "001110001",
11466 => "001100111",
11467 => "001100000",
11468 => "001100111",
11469 => "001101011",
11470 => "001110110",
11471 => "001101110",
11472 => "001101101",
11473 => "001110000",
11474 => "001101110",
11475 => "001100101",
11476 => "001100110",
11477 => "001101010",
11478 => "001101000",
11479 => "001101010",
11480 => "001111001",
11481 => "001111001",
11482 => "001110000",
11483 => "001110000",
11484 => "001110010",
11485 => "001110001",
11486 => "001110001",
11487 => "001110000",
11488 => "001100111",
11489 => "001110001",
11490 => "001110001",
11491 => "001110101",
11492 => "001110000",
11493 => "001100110",
11494 => "001011011",
11495 => "001100011",
11496 => "001100011",
11497 => "001100101",
11498 => "001011111",
11499 => "001010111",
11500 => "001011010",
11501 => "001011011",
11502 => "001011000",
11503 => "001011000",
11504 => "001100010",
11505 => "001011000",
11506 => "001011100",
11507 => "001010111",
11508 => "001011110",
11509 => "001011100",
11510 => "001011001",
11511 => "001010111",
11512 => "001010011",
11513 => "001010110",
11514 => "001010110",
11515 => "001011101",
11516 => "001011100",
11517 => "001011001",
11518 => "001010111",
11519 => "001011010",
11520 => "001000011",
11521 => "001001111",
11522 => "001000000",
11523 => "001001110",
11524 => "000110110",
11525 => "000111000",
11526 => "000101011",
11527 => "000110101",
11528 => "001000101",
11529 => "001000101",
11530 => "001100001",
11531 => "001100110",
11532 => "001001110",
11533 => "001001011",
11534 => "001001010",
11535 => "001001100",
11536 => "001001101",
11537 => "001100110",
11538 => "001100111",
11539 => "001011110",
11540 => "001101001",
11541 => "001100011",
11542 => "001011001",
11543 => "001010011",
11544 => "001000100",
11545 => "001001101",
11546 => "001011000",
11547 => "001011110",
11548 => "001011000",
11549 => "001011111",
11550 => "001011000",
11551 => "001100000",
11552 => "001101010",
11553 => "001100111",
11554 => "001100101",
11555 => "001101100",
11556 => "001100110",
11557 => "001100001",
11558 => "001011110",
11559 => "001010101",
11560 => "001011000",
11561 => "001010011",
11562 => "001010011",
11563 => "001101010",
11564 => "001100101",
11565 => "001011101",
11566 => "001100010",
11567 => "001100001",
11568 => "001100001",
11569 => "001100110",
11570 => "001101011",
11571 => "001101100",
11572 => "001101001",
11573 => "001101000",
11574 => "001100010",
11575 => "001100110",
11576 => "001011111",
11577 => "001101001",
11578 => "001011111",
11579 => "001011000",
11580 => "001100100",
11581 => "001100000",
11582 => "001100101",
11583 => "001100011",
11584 => "001011011",
11585 => "001100110",
11586 => "001101000",
11587 => "001101110",
11588 => "001101011",
11589 => "001101011",
11590 => "001101101",
11591 => "001110010",
11592 => "001100011",
11593 => "001101011",
11594 => "001101011",
11595 => "001101101",
11596 => "001100111",
11597 => "001101001",
11598 => "001101101",
11599 => "001100111",
11600 => "001101011",
11601 => "001101011",
11602 => "001100100",
11603 => "001100110",
11604 => "001100000",
11605 => "001101101",
11606 => "001101100",
11607 => "001101011",
11608 => "001101110",
11609 => "001101010",
11610 => "001101101",
11611 => "001101111",
11612 => "001110000",
11613 => "001101110",
11614 => "001101001",
11615 => "001101101",
11616 => "001100111",
11617 => "001100111",
11618 => "001101001",
11619 => "001101111",
11620 => "001100111",
11621 => "001101010",
11622 => "001101001",
11623 => "001100111",
11624 => "001100011",
11625 => "001101101",
11626 => "001011110",
11627 => "001011110",
11628 => "001011010",
11629 => "001011101",
11630 => "001100010",
11631 => "001011101",
11632 => "001100010",
11633 => "001100010",
11634 => "001100101",
11635 => "001010101",
11636 => "001011000",
11637 => "001010011",
11638 => "001011100",
11639 => "001011111",
11640 => "001010100",
11641 => "001010110",
11642 => "001001000",
11643 => "001011000",
11644 => "001001101",
11645 => "001000100",
11646 => "001010010",
11647 => "001001110",
11648 => "001001001",
11649 => "001010000",
11650 => "001011110",
11651 => "001000011",
11652 => "000110001",
11653 => "000101100",
11654 => "000101011",
11655 => "000100010",
11656 => "000110011",
11657 => "000101000",
11658 => "001010000",
11659 => "000110110",
11660 => "001001111",
11661 => "000111001",
11662 => "000110111",
11663 => "000110101",
11664 => "001010001",
11665 => "001110010",
11666 => "001110100",
11667 => "001100110",
11668 => "001100111",
11669 => "001100010",
11670 => "001100000",
11671 => "001100010",
11672 => "001100101",
11673 => "001100000",
11674 => "001011001",
11675 => "001100000",
11676 => "001011011",
11677 => "001010001",
11678 => "001011111",
11679 => "001011110",
11680 => "001010110",
11681 => "001011101",
11682 => "001011011",
11683 => "001011101",
11684 => "001100001",
11685 => "001100111",
11686 => "001100000",
11687 => "001011111",
11688 => "001101000",
11689 => "001101101",
11690 => "001010010",
11691 => "001010101",
11692 => "001001110",
11693 => "001011110",
11694 => "001011111",
11695 => "001011101",
11696 => "001100001",
11697 => "001011111",
11698 => "001100100",
11699 => "001101000",
11700 => "001100111",
11701 => "001100010",
11702 => "001011011",
11703 => "001101110",
11704 => "001011011",
11705 => "001100110",
11706 => "001100000",
11707 => "001100101",
11708 => "001101000",
11709 => "001100011",
11710 => "001100111",
11711 => "001101000",
11712 => "001101110",
11713 => "001100111",
11714 => "001101011",
11715 => "001100010",
11716 => "001100111",
11717 => "001100111",
11718 => "001100010",
11719 => "001110110",
11720 => "001101011",
11721 => "001100011",
11722 => "001100100",
11723 => "001100000",
11724 => "001100101",
11725 => "001100001",
11726 => "001100011",
11727 => "001101010",
11728 => "001100110",
11729 => "001100011",
11730 => "001101101",
11731 => "001100111",
11732 => "001110011",
11733 => "001101000",
11734 => "001101111",
11735 => "001011111",
11736 => "001011111",
11737 => "001101000",
11738 => "001100111",
11739 => "001101100",
11740 => "001100101",
11741 => "001100101",
11742 => "001101000",
11743 => "001101011",
11744 => "001101001",
11745 => "001100110",
11746 => "001011010",
11747 => "001010100",
11748 => "001011111",
11749 => "001100110",
11750 => "001100100",
11751 => "001100001",
11752 => "001101001",
11753 => "001101110",
11754 => "001101111",
11755 => "001101111",
11756 => "001100000",
11757 => "001100010",
11758 => "001011100",
11759 => "001011011",
11760 => "001010111",
11761 => "001011000",
11762 => "001011010",
11763 => "001100010",
11764 => "001011101",
11765 => "001100000",
11766 => "001011110",
11767 => "001010100",
11768 => "001010011",
11769 => "001010111",
11770 => "001001100",
11771 => "001001011",
11772 => "001010010",
11773 => "001000100",
11774 => "001001110",
11775 => "001001110",
11776 => "001010110",
11777 => "001011100",
11778 => "001011000",
11779 => "001001111",
11780 => "001010000",
11781 => "001001010",
11782 => "000111101",
11783 => "000011100",
11784 => "000111010",
11785 => "001000010",
11786 => "000110111",
11787 => "001001110",
11788 => "001001110",
11789 => "001001010",
11790 => "001001110",
11791 => "001010000",
11792 => "001011110",
11793 => "001101001",
11794 => "001111011",
11795 => "001101100",
11796 => "001101010",
11797 => "001100001",
11798 => "001100110",
11799 => "001101001",
11800 => "001101011",
11801 => "001101010",
11802 => "001100010",
11803 => "001100011",
11804 => "001011110",
11805 => "001100010",
11806 => "001100101",
11807 => "001100100",
11808 => "001011011",
11809 => "001100111",
11810 => "001011101",
11811 => "001010010",
11812 => "001010100",
11813 => "001011011",
11814 => "001100001",
11815 => "001100011",
11816 => "001100001",
11817 => "001100001",
11818 => "001101000",
11819 => "001010101",
11820 => "001010110",
11821 => "001010100",
11822 => "001010011",
11823 => "001011011",
11824 => "001010111",
11825 => "001011011",
11826 => "001011100",
11827 => "001011111",
11828 => "001011100",
11829 => "001100100",
11830 => "001100011",
11831 => "001100000",
11832 => "001100101",
11833 => "001100111",
11834 => "001100011",
11835 => "001101011",
11836 => "001110011",
11837 => "001101011",
11838 => "001101110",
11839 => "001110110",
11840 => "001101011",
11841 => "001110001",
11842 => "001101001",
11843 => "001100011",
11844 => "001101010",
11845 => "001100011",
11846 => "001100011",
11847 => "001101001",
11848 => "001110001",
11849 => "001100101",
11850 => "001100000",
11851 => "001011111",
11852 => "001100000",
11853 => "001011010",
11854 => "001100001",
11855 => "001011011",
11856 => "001100101",
11857 => "001100101",
11858 => "001011001",
11859 => "001011110",
11860 => "001100010",
11861 => "001100010",
11862 => "001101000",
11863 => "001100100",
11864 => "001011110",
11865 => "001011110",
11866 => "001100001",
11867 => "001011101",
11868 => "001011001",
11869 => "001101011",
11870 => "001101001",
11871 => "001100111",
11872 => "001101000",
11873 => "001100111",
11874 => "001100101",
11875 => "001101100",
11876 => "001101010",
11877 => "001100110",
11878 => "001100111",
11879 => "001100101",
11880 => "001100000",
11881 => "001101010",
11882 => "001011111",
11883 => "001101010",
11884 => "001100110",
11885 => "001101110",
11886 => "001100100",
11887 => "001011001",
11888 => "001011010",
11889 => "001011110",
11890 => "001011110",
11891 => "001010110",
11892 => "001100110",
11893 => "001100011",
11894 => "001011100",
11895 => "001011001",
11896 => "001011101",
11897 => "001011100",
11898 => "001011001",
11899 => "001010111",
11900 => "001010010",
11901 => "001011010",
11902 => "001011000",
11903 => "001010100",
11904 => "001011001",
11905 => "001011001",
11906 => "001100001",
11907 => "001001111",
11908 => "001001001",
11909 => "001001111",
11910 => "001001010",
11911 => "001010101",
11912 => "001010010",
11913 => "001010011",
11914 => "000111011",
11915 => "001000111",
11916 => "001010101",
11917 => "000100110",
11918 => "001001100",
11919 => "001000011",
11920 => "001100011",
11921 => "001011100",
11922 => "001101001",
11923 => "001110010",
11924 => "001011111",
11925 => "001011111",
11926 => "001110111",
11927 => "001100001",
11928 => "001100101",
11929 => "001011110",
11930 => "001100011",
11931 => "001100011",
11932 => "001011000",
11933 => "001011111",
11934 => "001011110",
11935 => "001011000",
11936 => "001001011",
11937 => "001010111",
11938 => "001010101",
11939 => "001011011",
11940 => "001100001",
11941 => "001011101",
11942 => "001011101",
11943 => "001011100",
11944 => "001011111",
11945 => "001100100",
11946 => "001100101",
11947 => "001101001",
11948 => "001101000",
11949 => "001110110",
11950 => "001100101",
11951 => "001100000",
11952 => "001100011",
11953 => "001100011",
11954 => "001100001",
11955 => "001010111",
11956 => "001100000",
11957 => "001011110",
11958 => "001010100",
11959 => "001011100",
11960 => "001011110",
11961 => "001101000",
11962 => "001101010",
11963 => "001100000",
11964 => "001011001",
11965 => "001100011",
11966 => "001100111",
11967 => "001100111",
11968 => "001101001",
11969 => "001100110",
11970 => "001100101",
11971 => "001101000",
11972 => "001100100",
11973 => "001100110",
11974 => "001100111",
11975 => "001101001",
11976 => "001101100",
11977 => "001100101",
11978 => "001011101",
11979 => "001010110",
11980 => "001100001",
11981 => "001011111",
11982 => "001011110",
11983 => "001011110",
11984 => "001011001",
11985 => "001011110",
11986 => "001010111",
11987 => "001010111",
11988 => "001011100",
11989 => "001011101",
11990 => "001010100",
11991 => "001011110",
11992 => "001011111",
11993 => "001011111",
11994 => "001100001",
11995 => "001100010",
11996 => "001100100",
11997 => "001011111",
11998 => "001100011",
11999 => "001100011",
12000 => "001100011",
12001 => "001101010",
12002 => "001100101",
12003 => "001100101",
12004 => "001100110",
12005 => "001100100",
12006 => "001101011",
12007 => "001101001",
12008 => "001100000",
12009 => "001101011",
12010 => "001101011",
12011 => "001100111",
12012 => "001101011",
12013 => "001100111",
12014 => "001101101",
12015 => "001011111",
12016 => "001011100",
12017 => "001101000",
12018 => "001101011",
12019 => "001101010",
12020 => "001100001",
12021 => "001011100",
12022 => "001011011",
12023 => "001011010",
12024 => "001001111",
12025 => "001011000",
12026 => "001100010",
12027 => "001010011",
12028 => "001001110",
12029 => "001010100",
12030 => "001010111",
12031 => "001000111",
12032 => "001010100",
12033 => "001011010",
12034 => "001011001",
12035 => "001011111",
12036 => "001010111",
12037 => "001001001",
12038 => "000111001",
12039 => "001001001",
12040 => "001001010",
12041 => "001010100",
12042 => "001011001",
12043 => "000011100",
12044 => "000100001",
12045 => "000110101",
12046 => "000101010",
12047 => "001011110",
12048 => "001100111",
12049 => "001110111",
12050 => "001101001",
12051 => "001011110",
12052 => "001101100",
12053 => "001100110",
12054 => "001111010",
12055 => "001011000",
12056 => "001101100",
12057 => "001101010",
12058 => "001100001",
12059 => "001100001",
12060 => "001011011",
12061 => "001011110",
12062 => "001010000",
12063 => "001000010",
12064 => "001001110",
12065 => "001010010",
12066 => "001100010",
12067 => "001100001",
12068 => "001011110",
12069 => "001011100",
12070 => "001010100",
12071 => "001100001",
12072 => "001100111",
12073 => "001101111",
12074 => "001101011",
12075 => "001100010",
12076 => "001100000",
12077 => "001100101",
12078 => "001100011",
12079 => "001010110",
12080 => "001001011",
12081 => "001100100",
12082 => "001100011",
12083 => "001101011",
12084 => "001100100",
12085 => "001100010",
12086 => "001011110",
12087 => "001100111",
12088 => "001011101",
12089 => "001011101",
12090 => "001100000",
12091 => "001100010",
12092 => "001101010",
12093 => "001101000",
12094 => "001100110",
12095 => "001101011",
12096 => "001101111",
12097 => "001100111",
12098 => "001100110",
12099 => "001100010",
12100 => "001100011",
12101 => "001101001",
12102 => "001100100",
12103 => "001100100",
12104 => "001100100",
12105 => "001100110",
12106 => "001100110",
12107 => "001011101",
12108 => "001010101",
12109 => "001011011",
12110 => "001100101",
12111 => "001100111",
12112 => "001011000",
12113 => "001010110",
12114 => "001100100",
12115 => "001011011",
12116 => "001001101",
12117 => "001010011",
12118 => "001011011",
12119 => "001100010",
12120 => "001011111",
12121 => "001011101",
12122 => "001011111",
12123 => "001011011",
12124 => "001010000",
12125 => "001100001",
12126 => "001011111",
12127 => "001100010",
12128 => "001100011",
12129 => "001011111",
12130 => "001100011",
12131 => "001011111",
12132 => "001100100",
12133 => "001100101",
12134 => "001100011",
12135 => "001100010",
12136 => "001100010",
12137 => "001100101",
12138 => "001011110",
12139 => "001011111",
12140 => "001100111",
12141 => "001011101",
12142 => "001010111",
12143 => "001100010",
12144 => "001100011",
12145 => "001100100",
12146 => "001011101",
12147 => "001011110",
12148 => "001100000",
12149 => "001100001",
12150 => "001100000",
12151 => "001100100",
12152 => "001100001",
12153 => "001011110",
12154 => "001010111",
12155 => "001100011",
12156 => "001011010",
12157 => "001010110",
12158 => "001011100",
12159 => "001010001",
12160 => "001011111",
12161 => "001101000",
12162 => "001010010",
12163 => "001011101",
12164 => "001101010",
12165 => "001010001",
12166 => "001011010",
12167 => "001001000",
12168 => "001001010",
12169 => "001000011",
12170 => "000100011",
12171 => "000101110",
12172 => "000100101",
12173 => "000101001",
12174 => "000110010",
12175 => "001010101",
12176 => "001001100",
12177 => "001111010",
12178 => "000111110",
12179 => "001011110",
12180 => "001010100",
12181 => "001011000",
12182 => "001111010",
12183 => "001100111",
12184 => "001101101",
12185 => "001100011",
12186 => "001010000",
12187 => "001100001",
12188 => "001011000",
12189 => "001010100",
12190 => "001011001",
12191 => "001010111",
12192 => "001011111",
12193 => "001100001",
12194 => "001011001",
12195 => "001100111",
12196 => "001100011",
12197 => "001011011",
12198 => "001010111",
12199 => "001100011",
12200 => "001100011",
12201 => "001011111",
12202 => "001011110",
12203 => "001101011",
12204 => "001011001",
12205 => "001100010",
12206 => "001100010",
12207 => "001100011",
12208 => "001101001",
12209 => "001100011",
12210 => "001100010",
12211 => "001100000",
12212 => "001100001",
12213 => "001100000",
12214 => "001010111",
12215 => "001011000",
12216 => "001011101",
12217 => "001101001",
12218 => "001100100",
12219 => "001101011",
12220 => "001011111",
12221 => "001100000",
12222 => "001100011",
12223 => "001100111",
12224 => "001101010",
12225 => "001100110",
12226 => "001011101",
12227 => "001101011",
12228 => "001100101",
12229 => "001100100",
12230 => "001101011",
12231 => "001101010",
12232 => "001101100",
12233 => "001101010",
12234 => "001101010",
12235 => "001101010",
12236 => "001100111",
12237 => "001100101",
12238 => "001100010",
12239 => "001100101",
12240 => "001100110",
12241 => "001100101",
12242 => "001101000",
12243 => "001100010",
12244 => "001100010",
12245 => "001100110",
12246 => "001100100",
12247 => "001100101",
12248 => "001100000",
12249 => "001011100",
12250 => "001010101",
12251 => "001011100",
12252 => "001011010",
12253 => "001100001",
12254 => "001100000",
12255 => "001100010",
12256 => "001011111",
12257 => "001011010",
12258 => "001011010",
12259 => "001011010",
12260 => "001011100",
12261 => "001100001",
12262 => "001011010",
12263 => "001010100",
12264 => "001011100",
12265 => "001011100",
12266 => "001100100",
12267 => "001011110",
12268 => "001011110",
12269 => "001100110",
12270 => "001100001",
12271 => "001100100",
12272 => "001011100",
12273 => "001011100",
12274 => "001100100",
12275 => "001100100",
12276 => "001101000",
12277 => "001100000",
12278 => "001100110",
12279 => "001100111",
12280 => "001100001",
12281 => "001100000",
12282 => "001100000",
12283 => "001011000",
12284 => "001011010",
12285 => "001011000",
12286 => "001011000",
12287 => "001011010",
12288 => "001100010",
12289 => "001101001",
12290 => "001011010",
12291 => "001100110",
12292 => "001011110",
12293 => "001010110",
12294 => "001101001",
12295 => "001011000",
12296 => "001001111",
12297 => "000110011",
12298 => "000110101",
12299 => "001000001",
12300 => "000110001",
12301 => "000101100",
12302 => "000110110",
12303 => "000110110",
12304 => "001100100",
12305 => "001100010",
12306 => "001001101",
12307 => "001100000",
12308 => "001101010",
12309 => "001110010",
12310 => "001001000",
12311 => "001001011",
12312 => "001100000",
12313 => "001011000",
12314 => "001101000",
12315 => "001011010",
12316 => "001011111",
12317 => "001010100",
12318 => "001010110",
12319 => "001011010",
12320 => "001101010",
12321 => "001100110",
12322 => "001100101",
12323 => "001100110",
12324 => "001100110",
12325 => "001011010",
12326 => "001011001",
12327 => "001011001",
12328 => "001011001",
12329 => "001010100",
12330 => "001011101",
12331 => "001010010",
12332 => "001010110",
12333 => "001100000",
12334 => "001100100",
12335 => "001011100",
12336 => "001100100",
12337 => "001100110",
12338 => "001100011",
12339 => "001011100",
12340 => "001011101",
12341 => "001101010",
12342 => "001100110",
12343 => "001011100",
12344 => "001011000",
12345 => "001011001",
12346 => "001011101",
12347 => "001101001",
12348 => "001101010",
12349 => "001100010",
12350 => "001100000",
12351 => "001101010",
12352 => "001101100",
12353 => "001101010",
12354 => "001110010",
12355 => "001101010",
12356 => "001100010",
12357 => "001010101",
12358 => "001011111",
12359 => "001110110",
12360 => "001101001",
12361 => "001101000",
12362 => "001011001",
12363 => "001011100",
12364 => "001011010",
12365 => "001011111",
12366 => "001011111",
12367 => "001011010",
12368 => "001100000",
12369 => "001011011",
12370 => "001011001",
12371 => "001011100",
12372 => "001100101",
12373 => "001100010",
12374 => "001100111",
12375 => "001100101",
12376 => "001100010",
12377 => "001100100",
12378 => "001100100",
12379 => "001100010",
12380 => "001100101",
12381 => "001100001",
12382 => "001101001",
12383 => "001100000",
12384 => "001011110",
12385 => "001100010",
12386 => "001100011",
12387 => "001011101",
12388 => "001001101",
12389 => "001001100",
12390 => "001010010",
12391 => "001010110",
12392 => "001011110",
12393 => "001011100",
12394 => "001011010",
12395 => "001100000",
12396 => "001011101",
12397 => "001011001",
12398 => "001011101",
12399 => "001011101",
12400 => "001100000",
12401 => "001010001",
12402 => "001011011",
12403 => "001100100",
12404 => "001101000",
12405 => "001100100",
12406 => "001100000",
12407 => "001101001",
12408 => "001101011",
12409 => "001100100",
12410 => "001100010",
12411 => "001100100",
12412 => "001100110",
12413 => "001011000",
12414 => "001011110",
12415 => "001001001",
12416 => "001011010",
12417 => "001011111",
12418 => "001100100",
12419 => "001011100",
12420 => "001011110",
12421 => "001011101",
12422 => "001100000",
12423 => "001010111",
12424 => "001010100",
12425 => "001010000",
12426 => "000111111",
12427 => "000110010",
12428 => "000111100",
12429 => "000100101",
12430 => "000101010",
12431 => "000101100",
12432 => "001100100",
12433 => "001010111",
12434 => "001011000",
12435 => "001011000",
12436 => "001011100",
12437 => "001100101",
12438 => "001100101",
12439 => "001010101",
12440 => "001000011",
12441 => "001100100",
12442 => "001100100",
12443 => "001100111",
12444 => "001100011",
12445 => "001101011",
12446 => "001110100",
12447 => "001111111",
12448 => "001110101",
12449 => "001100111",
12450 => "001101110",
12451 => "001011101",
12452 => "001101000",
12453 => "001100100",
12454 => "001100011",
12455 => "001011111",
12456 => "001100001",
12457 => "001100100",
12458 => "010000000",
12459 => "001011110",
12460 => "001100001",
12461 => "001101000",
12462 => "001100001",
12463 => "001100101",
12464 => "001011110",
12465 => "001011011",
12466 => "001100010",
12467 => "001100100",
12468 => "001100010",
12469 => "001100101",
12470 => "001100111",
12471 => "001101100",
12472 => "001101010",
12473 => "001100101",
12474 => "001011000",
12475 => "001011011",
12476 => "001011001",
12477 => "001011011",
12478 => "001100010",
12479 => "001010110",
12480 => "001010110",
12481 => "001011100",
12482 => "001100100",
12483 => "001100101",
12484 => "001101111",
12485 => "001101000",
12486 => "001100111",
12487 => "001100110",
12488 => "001100001",
12489 => "001011010",
12490 => "001011010",
12491 => "001011101",
12492 => "001100001",
12493 => "001100011",
12494 => "001010110",
12495 => "001010010",
12496 => "001100000",
12497 => "001011110",
12498 => "001011010",
12499 => "001100010",
12500 => "001100101",
12501 => "001100110",
12502 => "001100100",
12503 => "001100011",
12504 => "001100000",
12505 => "001100100",
12506 => "001101010",
12507 => "001100100",
12508 => "001100000",
12509 => "001011111",
12510 => "001100000",
12511 => "001011101",
12512 => "001011011",
12513 => "001011001",
12514 => "001100100",
12515 => "001101000",
12516 => "001011101",
12517 => "001010110",
12518 => "001010010",
12519 => "001001011",
12520 => "001010110",
12521 => "001010101",
12522 => "001001111",
12523 => "001011100",
12524 => "001100001",
12525 => "001011101",
12526 => "001011100",
12527 => "001011101",
12528 => "001011101",
12529 => "001100100",
12530 => "001011101",
12531 => "001011101",
12532 => "001011001",
12533 => "001100000",
12534 => "001011101",
12535 => "001011011",
12536 => "001010001",
12537 => "001011001",
12538 => "001011101",
12539 => "001100010",
12540 => "001011110",
12541 => "001100010",
12542 => "001100011",
12543 => "001100000",
12544 => "001010110",
12545 => "001010111",
12546 => "001010101",
12547 => "001011011",
12548 => "001100010",
12549 => "001011011",
12550 => "001011111",
12551 => "001011111",
12552 => "001011100",
12553 => "001011010",
12554 => "001010110",
12555 => "001010100",
12556 => "001001100",
12557 => "001001001",
12558 => "000111110",
12559 => "000110110",
12560 => "001100100",
12561 => "001011001",
12562 => "000111011",
12563 => "001000111",
12564 => "000110111",
12565 => "001001000",
12566 => "001001101",
12567 => "000101001",
12568 => "001000101",
12569 => "000011111",
12570 => "001000011",
12571 => "001010100",
12572 => "001101111",
12573 => "001100001",
12574 => "001111111",
12575 => "001111000",
12576 => "001100000",
12577 => "010000111",
12578 => "001011111",
12579 => "001111111",
12580 => "001100000",
12581 => "001101000",
12582 => "001011101",
12583 => "001100000",
12584 => "001011101",
12585 => "001100011",
12586 => "001111001",
12587 => "001101101",
12588 => "001100101",
12589 => "001100011",
12590 => "001010000",
12591 => "001010100",
12592 => "001101000",
12593 => "001100011",
12594 => "001011001",
12595 => "001011000",
12596 => "001011111",
12597 => "001100011",
12598 => "001011111",
12599 => "001100011",
12600 => "001011011",
12601 => "001101001",
12602 => "001101000",
12603 => "001101101",
12604 => "001100111",
12605 => "001100001",
12606 => "001011110",
12607 => "001100100",
12608 => "001100001",
12609 => "001011011",
12610 => "001100101",
12611 => "001101000",
12612 => "001101010",
12613 => "001100001",
12614 => "001100010",
12615 => "001011101",
12616 => "001100001",
12617 => "001011111",
12618 => "001011110",
12619 => "001011101",
12620 => "001011111",
12621 => "001100000",
12622 => "001100100",
12623 => "001011010",
12624 => "001010101",
12625 => "001011011",
12626 => "001011110",
12627 => "001011000",
12628 => "001010111",
12629 => "001011001",
12630 => "001011000",
12631 => "001100010",
12632 => "001101000",
12633 => "001100101",
12634 => "001100010",
12635 => "001100110",
12636 => "001100011",
12637 => "001100010",
12638 => "001100010",
12639 => "001100001",
12640 => "001011111",
12641 => "001011000",
12642 => "001010110",
12643 => "001011101",
12644 => "001100000",
12645 => "001100001",
12646 => "001010100",
12647 => "001010111",
12648 => "001010110",
12649 => "001011110",
12650 => "001011000",
12651 => "001010001",
12652 => "001010001",
12653 => "001011011",
12654 => "001011110",
12655 => "001100100",
12656 => "001011100",
12657 => "001010111",
12658 => "001011001",
12659 => "001011011",
12660 => "001011101",
12661 => "001011110",
12662 => "001100000",
12663 => "001010011",
12664 => "001011100",
12665 => "001011010",
12666 => "001011001",
12667 => "001011001",
12668 => "001011101",
12669 => "001100000",
12670 => "001011011",
12671 => "001011010",
12672 => "001010110",
12673 => "001011000",
12674 => "001010100",
12675 => "001010111",
12676 => "001011101",
12677 => "001010111",
12678 => "001011000",
12679 => "001100010",
12680 => "001100000",
12681 => "001100100",
12682 => "001010100",
12683 => "001010101",
12684 => "001010111",
12685 => "001011101",
12686 => "000111000",
12687 => "001000110",
12688 => "001101011",
12689 => "001000011",
12690 => "000110001",
12691 => "001001010",
12692 => "001000101",
12693 => "001000001",
12694 => "000110100",
12695 => "000111000",
12696 => "001100001",
12697 => "001110110",
12698 => "000110101",
12699 => "001000111",
12700 => "001100010",
12701 => "001100110",
12702 => "001100101",
12703 => "001110000",
12704 => "001001001",
12705 => "000111000",
12706 => "001101100",
12707 => "001101100",
12708 => "001101101",
12709 => "001101111",
12710 => "001101111",
12711 => "001100110",
12712 => "001100101",
12713 => "001100000",
12714 => "001100100",
12715 => "001100000",
12716 => "001011001",
12717 => "001100011",
12718 => "001110101",
12719 => "001011001",
12720 => "001011100",
12721 => "001100100",
12722 => "001101011",
12723 => "001101000",
12724 => "001101000",
12725 => "001101001",
12726 => "001100110",
12727 => "001100100",
12728 => "001100101",
12729 => "001100111",
12730 => "001100011",
12731 => "001100011",
12732 => "001101010",
12733 => "001101000",
12734 => "001101000",
12735 => "001101100",
12736 => "001100110",
12737 => "001101001",
12738 => "001101010",
12739 => "001011010",
12740 => "001100011",
12741 => "001100011",
12742 => "001100100",
12743 => "001100101",
12744 => "001101001",
12745 => "001100100",
12746 => "001011111",
12747 => "001100100",
12748 => "001011111",
12749 => "001010101",
12750 => "001001101",
12751 => "001100011",
12752 => "001101011",
12753 => "001100101",
12754 => "001100110",
12755 => "001101010",
12756 => "001100110",
12757 => "001010101",
12758 => "001010000",
12759 => "001000001",
12760 => "001010000",
12761 => "001011110",
12762 => "001100011",
12763 => "001011111",
12764 => "001100001",
12765 => "001100111",
12766 => "001100011",
12767 => "001100100",
12768 => "001100000",
12769 => "001011101",
12770 => "001011110",
12771 => "001011101",
12772 => "001011000",
12773 => "001011011",
12774 => "001011001",
12775 => "001011010",
12776 => "001011011",
12777 => "001011100",
12778 => "001100001",
12779 => "001011010",
12780 => "001001111",
12781 => "001010001",
12782 => "001010101",
12783 => "001011010",
12784 => "001011010",
12785 => "001011000",
12786 => "001010100",
12787 => "001011001",
12788 => "001010011",
12789 => "001010111",
12790 => "001100000",
12791 => "001011110",
12792 => "001100010",
12793 => "001011110",
12794 => "001010100",
12795 => "001010011",
12796 => "001100011",
12797 => "001100010",
12798 => "001010110",
12799 => "001011011",
12800 => "001010100",
12801 => "001100011",
12802 => "001001010",
12803 => "001010100",
12804 => "001010011",
12805 => "001011001",
12806 => "001011011",
12807 => "001101001",
12808 => "001100000",
12809 => "001100100",
12810 => "001100100",
12811 => "001100001",
12812 => "001100101",
12813 => "001101000",
12814 => "001100110",
12815 => "001100100",
12816 => "001011001",
12817 => "001100001",
12818 => "001001010",
12819 => "001010000",
12820 => "001010011",
12821 => "001010100",
12822 => "001011111",
12823 => "000111110",
12824 => "010001100",
12825 => "001101001",
12826 => "010000101",
12827 => "000111101",
12828 => "001010011",
12829 => "001010001",
12830 => "001010011",
12831 => "001101010",
12832 => "001001011",
12833 => "001101101",
12834 => "001111011",
12835 => "001100010",
12836 => "010001001",
12837 => "001110100",
12838 => "010000010",
12839 => "001100110",
12840 => "001011011",
12841 => "001100110",
12842 => "001110100",
12843 => "001011110",
12844 => "001011101",
12845 => "001010011",
12846 => "001101110",
12847 => "001100111",
12848 => "001101101",
12849 => "001100011",
12850 => "001100110",
12851 => "001100111",
12852 => "001011111",
12853 => "001100101",
12854 => "001100000",
12855 => "001100001",
12856 => "001100100",
12857 => "001101011",
12858 => "001100010",
12859 => "001100101",
12860 => "001100101",
12861 => "001100010",
12862 => "001100101",
12863 => "001011100",
12864 => "001101101",
12865 => "001101100",
12866 => "001100110",
12867 => "001100011",
12868 => "001011011",
12869 => "001100010",
12870 => "001011111",
12871 => "001101010",
12872 => "001101001",
12873 => "001101111",
12874 => "001101001",
12875 => "001100111",
12876 => "001100110",
12877 => "001100110",
12878 => "001100010",
12879 => "001101010",
12880 => "001101111",
12881 => "001100011",
12882 => "001101001",
12883 => "001101001",
12884 => "001101001",
12885 => "001011111",
12886 => "001100000",
12887 => "001011101",
12888 => "001011011",
12889 => "001100000",
12890 => "001100101",
12891 => "001100011",
12892 => "001011011",
12893 => "001011101",
12894 => "001011011",
12895 => "001011010",
12896 => "001011101",
12897 => "001011100",
12898 => "001100010",
12899 => "001100000",
12900 => "001011100",
12901 => "001011110",
12902 => "001001110",
12903 => "001010111",
12904 => "001010111",
12905 => "001100000",
12906 => "001100010",
12907 => "001100110",
12908 => "001100100",
12909 => "001011100",
12910 => "001011010",
12911 => "001011000",
12912 => "001011101",
12913 => "001100001",
12914 => "001011010",
12915 => "001011100",
12916 => "001010011",
12917 => "001010110",
12918 => "001010011",
12919 => "001010110",
12920 => "001011010",
12921 => "001011000",
12922 => "001010010",
12923 => "001010011",
12924 => "001011100",
12925 => "001100100",
12926 => "001011010",
12927 => "001010111",
12928 => "001110001",
12929 => "001011100",
12930 => "001010110",
12931 => "001011010",
12932 => "001011100",
12933 => "001001100",
12934 => "001000100",
12935 => "001001111",
12936 => "001011101",
12937 => "001011111",
12938 => "001011101",
12939 => "001100111",
12940 => "001010001",
12941 => "001101011",
12942 => "001100110",
12943 => "001101110",
12944 => "001100100",
12945 => "001101101",
12946 => "001100111",
12947 => "001100010",
12948 => "001010101",
12949 => "001010101",
12950 => "001010000",
12951 => "001100111",
12952 => "010000010",
12953 => "001011101",
12954 => "001100010",
12955 => "001101101",
12956 => "001011111",
12957 => "001011010",
12958 => "001100011",
12959 => "001110101",
12960 => "001101101",
12961 => "001101111",
12962 => "001010010",
12963 => "001110010",
12964 => "010001000",
12965 => "010000001",
12966 => "010000001",
12967 => "010011010",
12968 => "001110010",
12969 => "010000000",
12970 => "001010101",
12971 => "001011011",
12972 => "010001110",
12973 => "010010110",
12974 => "001100001",
12975 => "001101101",
12976 => "001110011",
12977 => "001001111",
12978 => "001100010",
12979 => "001101110",
12980 => "001011101",
12981 => "001011110",
12982 => "001011111",
12983 => "001110010",
12984 => "001101111",
12985 => "001101011",
12986 => "001100001",
12987 => "001100011",
12988 => "001100001",
12989 => "001100001",
12990 => "001100000",
12991 => "001011011",
12992 => "001100110",
12993 => "001101000",
12994 => "001101001",
12995 => "001101001",
12996 => "001101010",
12997 => "001100010",
12998 => "001100110",
12999 => "001100111",
13000 => "001101101",
13001 => "001101010",
13002 => "001101011",
13003 => "001101101",
13004 => "001100110",
13005 => "001100100",
13006 => "001011101",
13007 => "001100011",
13008 => "001011010",
13009 => "001101000",
13010 => "001101000",
13011 => "001101010",
13012 => "001100110",
13013 => "001100001",
13014 => "001100111",
13015 => "001101000",
13016 => "001100101",
13017 => "001100000",
13018 => "001011101",
13019 => "001011111",
13020 => "001100010",
13021 => "001100000",
13022 => "001100010",
13023 => "001101100",
13024 => "001100100",
13025 => "001100010",
13026 => "001011110",
13027 => "001010110",
13028 => "001011001",
13029 => "001011100",
13030 => "001100101",
13031 => "001011110",
13032 => "001011100",
13033 => "001100000",
13034 => "001011110",
13035 => "001100000",
13036 => "001100110",
13037 => "001011100",
13038 => "001011100",
13039 => "001010101",
13040 => "001010111",
13041 => "001011011",
13042 => "001011110",
13043 => "001011011",
13044 => "001010110",
13045 => "001011011",
13046 => "001011011",
13047 => "001100000",
13048 => "001011001",
13049 => "001011101",
13050 => "001011101",
13051 => "001011110",
13052 => "001100001",
13053 => "001101011",
13054 => "001011111",
13055 => "001011000",
13056 => "001100110",
13057 => "001100101",
13058 => "001011111",
13059 => "001001000",
13060 => "001100101",
13061 => "001011010",
13062 => "001000110",
13063 => "001011000",
13064 => "001001100",
13065 => "001010000",
13066 => "001010010",
13067 => "001011101",
13068 => "001010100",
13069 => "001011000",
13070 => "001101011",
13071 => "001101101",
13072 => "001100011",
13073 => "001100100",
13074 => "001100011",
13075 => "001100011",
13076 => "001100000",
13077 => "001100011",
13078 => "001011111",
13079 => "001110100",
13080 => "010001000",
13081 => "001100111",
13082 => "000110111",
13083 => "001000000",
13084 => "001001011",
13085 => "001100101",
13086 => "001010000",
13087 => "001010101",
13088 => "010001110",
13089 => "001101101",
13090 => "001100000",
13091 => "010000000",
13092 => "001110100",
13093 => "001111001",
13094 => "001100111",
13095 => "001111010",
13096 => "001010101",
13097 => "001100011",
13098 => "001101110",
13099 => "000111010",
13100 => "001001001",
13101 => "001000111",
13102 => "010000101",
13103 => "001101100",
13104 => "010000010",
13105 => "010010010",
13106 => "010000101",
13107 => "010000111",
13108 => "001100110",
13109 => "001010010",
13110 => "001101000",
13111 => "001100100",
13112 => "001011110",
13113 => "001100100",
13114 => "001101000",
13115 => "001100001",
13116 => "001101000",
13117 => "001101001",
13118 => "001101011",
13119 => "001101111",
13120 => "001101001",
13121 => "001100011",
13122 => "001100100",
13123 => "001100010",
13124 => "001101011",
13125 => "001101001",
13126 => "001100011",
13127 => "001100100",
13128 => "001011110",
13129 => "001011101",
13130 => "001011110",
13131 => "001100100",
13132 => "001100101",
13133 => "001011101",
13134 => "001001010",
13135 => "001001101",
13136 => "001100100",
13137 => "001101011",
13138 => "001100111",
13139 => "001100010",
13140 => "001100010",
13141 => "001100110",
13142 => "001011100",
13143 => "001100000",
13144 => "001100001",
13145 => "001100011",
13146 => "001011110",
13147 => "001011111",
13148 => "001100001",
13149 => "001011101",
13150 => "001100010",
13151 => "001100110",
13152 => "001100001",
13153 => "001100010",
13154 => "001100000",
13155 => "001100110",
13156 => "001010111",
13157 => "001010100",
13158 => "001001000",
13159 => "001011110",
13160 => "001011011",
13161 => "001011001",
13162 => "001010111",
13163 => "001011000",
13164 => "001011101",
13165 => "001100010",
13166 => "001100100",
13167 => "001100001",
13168 => "001100001",
13169 => "001011101",
13170 => "001010010",
13171 => "001011011",
13172 => "001011010",
13173 => "001010101",
13174 => "001011001",
13175 => "001011111",
13176 => "001100000",
13177 => "001011101",
13178 => "001011110",
13179 => "001010011",
13180 => "001010100",
13181 => "001011010",
13182 => "001011010",
13183 => "001011110",
13184 => "001101001",
13185 => "001101100",
13186 => "001100100",
13187 => "001010101",
13188 => "001011001",
13189 => "001100100",
13190 => "001010001",
13191 => "001011001",
13192 => "001010110",
13193 => "001001011",
13194 => "001001001",
13195 => "001001110",
13196 => "001001111",
13197 => "001010010",
13198 => "001001000",
13199 => "001101101",
13200 => "001011001",
13201 => "001011100",
13202 => "001100000",
13203 => "001100100",
13204 => "001101001",
13205 => "001011001",
13206 => "001011001",
13207 => "001100101",
13208 => "001101101",
13209 => "001100001",
13210 => "001011100",
13211 => "001001110",
13212 => "001000001",
13213 => "001001101",
13214 => "001000110",
13215 => "001101011",
13216 => "010001011",
13217 => "010001101",
13218 => "010011100",
13219 => "001101001",
13220 => "001001101",
13221 => "010000001",
13222 => "001000000",
13223 => "001101010",
13224 => "010000111",
13225 => "001100001",
13226 => "000110111",
13227 => "001100101",
13228 => "001110101",
13229 => "001011111",
13230 => "001100000",
13231 => "001001010",
13232 => "001101011",
13233 => "010001000",
13234 => "001101110",
13235 => "001110001",
13236 => "001001110",
13237 => "001100111",
13238 => "001101010",
13239 => "001100111",
13240 => "001101000",
13241 => "001101010",
13242 => "001100100",
13243 => "001101010",
13244 => "001011110",
13245 => "001100101",
13246 => "001100110",
13247 => "001101010",
13248 => "001100111",
13249 => "001101001",
13250 => "001101010",
13251 => "001101101",
13252 => "001100100",
13253 => "001100010",
13254 => "001101011",
13255 => "001100000",
13256 => "001100000",
13257 => "001011001",
13258 => "001100000",
13259 => "001100001",
13260 => "001100101",
13261 => "001100100",
13262 => "001011100",
13263 => "001010100",
13264 => "001100011",
13265 => "001101010",
13266 => "001101011",
13267 => "001101101",
13268 => "001100111",
13269 => "001100011",
13270 => "001100010",
13271 => "001011111",
13272 => "001011100",
13273 => "001011011",
13274 => "001100001",
13275 => "001100001",
13276 => "001010101",
13277 => "001011010",
13278 => "001011110",
13279 => "001100101",
13280 => "001011110",
13281 => "001011101",
13282 => "001000111",
13283 => "001011101",
13284 => "001100101",
13285 => "001100000",
13286 => "001011100",
13287 => "001100110",
13288 => "001100000",
13289 => "001011110",
13290 => "001011110",
13291 => "001010100",
13292 => "001010100",
13293 => "001010011",
13294 => "001001101",
13295 => "001000110",
13296 => "001000110",
13297 => "001011011",
13298 => "001011010",
13299 => "001011110",
13300 => "001011010",
13301 => "001011001",
13302 => "001010011",
13303 => "001001110",
13304 => "001011010",
13305 => "001011101",
13306 => "001011100",
13307 => "001011001",
13308 => "001010100",
13309 => "001011110",
13310 => "001011000",
13311 => "001011010",
13312 => "001100111",
13313 => "001100111",
13314 => "001010011",
13315 => "001001011",
13316 => "001011011",
13317 => "001011100",
13318 => "001001100",
13319 => "001010000",
13320 => "001000001",
13321 => "001001111",
13322 => "001000100",
13323 => "001000101",
13324 => "001000110",
13325 => "000111111",
13326 => "001010011",
13327 => "001001011",
13328 => "001011100",
13329 => "001011111",
13330 => "001010010",
13331 => "001011111",
13332 => "001100001",
13333 => "001101000",
13334 => "001011101",
13335 => "001011011",
13336 => "001100110",
13337 => "001010111",
13338 => "001100000",
13339 => "001101001",
13340 => "001100110",
13341 => "001011010",
13342 => "010001011",
13343 => "001101101",
13344 => "001101100",
13345 => "001101011",
13346 => "001000110",
13347 => "001001000",
13348 => "001110011",
13349 => "001011110",
13350 => "001000111",
13351 => "000110011",
13352 => "001001101",
13353 => "001101000",
13354 => "001110011",
13355 => "010000010",
13356 => "001111010",
13357 => "010010000",
13358 => "001011111",
13359 => "001001011",
13360 => "001011001",
13361 => "001111111",
13362 => "001101110",
13363 => "001001010",
13364 => "010000000",
13365 => "001110111",
13366 => "001101011",
13367 => "001100101",
13368 => "001011010",
13369 => "001011000",
13370 => "001011111",
13371 => "001100011",
13372 => "001101011",
13373 => "001100110",
13374 => "001100101",
13375 => "001100010",
13376 => "001101100",
13377 => "001101011",
13378 => "001101001",
13379 => "001100101",
13380 => "001100111",
13381 => "001101001",
13382 => "001101000",
13383 => "001101000",
13384 => "001100100",
13385 => "001100001",
13386 => "001010010",
13387 => "001011101",
13388 => "001011001",
13389 => "001100000",
13390 => "001011100",
13391 => "001010111",
13392 => "001010111",
13393 => "001011111",
13394 => "001100000",
13395 => "001011100",
13396 => "001101010",
13397 => "001101010",
13398 => "001010110",
13399 => "001010011",
13400 => "001001000",
13401 => "001001111",
13402 => "001010101",
13403 => "001100000",
13404 => "001100010",
13405 => "001011011",
13406 => "001100111",
13407 => "001011011",
13408 => "001100001",
13409 => "001011111",
13410 => "001011111",
13411 => "001011100",
13412 => "001011111",
13413 => "001100110",
13414 => "001011011",
13415 => "001010100",
13416 => "001010011",
13417 => "001011010",
13418 => "001100110",
13419 => "001100000",
13420 => "001011101",
13421 => "001100010",
13422 => "001010111",
13423 => "001001101",
13424 => "001000110",
13425 => "001001010",
13426 => "001010001",
13427 => "001010000",
13428 => "001001111",
13429 => "001001110",
13430 => "001010010",
13431 => "001010101",
13432 => "001010010",
13433 => "001010100",
13434 => "001011110",
13435 => "001010011",
13436 => "001010101",
13437 => "001011001",
13438 => "001011011",
13439 => "001010110",
13440 => "001011010",
13441 => "001011011",
13442 => "001010101",
13443 => "001000101",
13444 => "001100000",
13445 => "001011000",
13446 => "001010001",
13447 => "001000101",
13448 => "000111000",
13449 => "000111010",
13450 => "001000000",
13451 => "000111100",
13452 => "000111111",
13453 => "001010100",
13454 => "001001001",
13455 => "001011001",
13456 => "001100010",
13457 => "001101010",
13458 => "001010101",
13459 => "001010011",
13460 => "001010101",
13461 => "001011110",
13462 => "001100111",
13463 => "001100101",
13464 => "001100110",
13465 => "001100000",
13466 => "001101010",
13467 => "001101010",
13468 => "001011011",
13469 => "001100111",
13470 => "001110000",
13471 => "001011101",
13472 => "000111111",
13473 => "000111010",
13474 => "001011110",
13475 => "001001110",
13476 => "001100100",
13477 => "001110100",
13478 => "000111100",
13479 => "001001010",
13480 => "000110011",
13481 => "001101000",
13482 => "001111000",
13483 => "001111100",
13484 => "001011011",
13485 => "001001011",
13486 => "001010001",
13487 => "000101101",
13488 => "000111111",
13489 => "001001001",
13490 => "001100000",
13491 => "010010011",
13492 => "000110111",
13493 => "010001011",
13494 => "001011111",
13495 => "001011001",
13496 => "001011100",
13497 => "001100000",
13498 => "001100001",
13499 => "001100101",
13500 => "001011111",
13501 => "001001100",
13502 => "000111101",
13503 => "001001110",
13504 => "001100110",
13505 => "001100010",
13506 => "001011011",
13507 => "001101000",
13508 => "001100110",
13509 => "001011111",
13510 => "001010101",
13511 => "001011101",
13512 => "001100000",
13513 => "001100101",
13514 => "001100110",
13515 => "001100000",
13516 => "001100000",
13517 => "001011110",
13518 => "001100100",
13519 => "001100010",
13520 => "001011111",
13521 => "001011011",
13522 => "001011010",
13523 => "001001110",
13524 => "001011010",
13525 => "001011111",
13526 => "001100010",
13527 => "001100011",
13528 => "001100011",
13529 => "001010110",
13530 => "001001010",
13531 => "001010000",
13532 => "001011001",
13533 => "001011101",
13534 => "001011011",
13535 => "001011011",
13536 => "001010100",
13537 => "001010011",
13538 => "001011010",
13539 => "001010100",
13540 => "001010001",
13541 => "001011100",
13542 => "001100011",
13543 => "001011110",
13544 => "001011000",
13545 => "001010001",
13546 => "001011001",
13547 => "001011100",
13548 => "001011011",
13549 => "001011100",
13550 => "001010000",
13551 => "001011010",
13552 => "001011010",
13553 => "001011011",
13554 => "001011110",
13555 => "001010101",
13556 => "001001110",
13557 => "001010010",
13558 => "001001110",
13559 => "001010011",
13560 => "001011010",
13561 => "001010110",
13562 => "001010011",
13563 => "001011010",
13564 => "001001101",
13565 => "001001111",
13566 => "001011000",
13567 => "001001111",
13568 => "001100000",
13569 => "001010010",
13570 => "001011001",
13571 => "001010001",
13572 => "001001100",
13573 => "001011010",
13574 => "001001100",
13575 => "001001000",
13576 => "000111101",
13577 => "000111110",
13578 => "000111010",
13579 => "000111000",
13580 => "000111010",
13581 => "001010010",
13582 => "001000111",
13583 => "001010111",
13584 => "001100010",
13585 => "001011100",
13586 => "001010101",
13587 => "001001101",
13588 => "001001101",
13589 => "001001011",
13590 => "001011001",
13591 => "001100001",
13592 => "001100001",
13593 => "001100000",
13594 => "001100100",
13595 => "001101111",
13596 => "001101100",
13597 => "001101100",
13598 => "001110000",
13599 => "001011100",
13600 => "001001111",
13601 => "000101000",
13602 => "001000001",
13603 => "001000111",
13604 => "000111000",
13605 => "001001001",
13606 => "000111111",
13607 => "001001110",
13608 => "000101110",
13609 => "001101110",
13610 => "001011110",
13611 => "000111011",
13612 => "001001101",
13613 => "000100011",
13614 => "001001010",
13615 => "001001000",
13616 => "001011001",
13617 => "001000000",
13618 => "001000110",
13619 => "001001011",
13620 => "001001110",
13621 => "000110111",
13622 => "001001001",
13623 => "001101110",
13624 => "001011010",
13625 => "001100111",
13626 => "001100000",
13627 => "001011100",
13628 => "001100111",
13629 => "001100001",
13630 => "001100010",
13631 => "001011100",
13632 => "001000000",
13633 => "001101110",
13634 => "001100100",
13635 => "001100011",
13636 => "001100001",
13637 => "001101100",
13638 => "001011100",
13639 => "001011001",
13640 => "001011000",
13641 => "001010011",
13642 => "001010111",
13643 => "001011111",
13644 => "001100001",
13645 => "001010011",
13646 => "001010010",
13647 => "001011010",
13648 => "001010010",
13649 => "001100101",
13650 => "001100111",
13651 => "001011111",
13652 => "001001001",
13653 => "001011000",
13654 => "001011100",
13655 => "001011010",
13656 => "001011110",
13657 => "001100011",
13658 => "001010111",
13659 => "001001001",
13660 => "001010110",
13661 => "001010101",
13662 => "001011011",
13663 => "001011101",
13664 => "001011000",
13665 => "001001100",
13666 => "001001100",
13667 => "001001011",
13668 => "001010101",
13669 => "001100111",
13670 => "001100100",
13671 => "001011111",
13672 => "001011110",
13673 => "001010100",
13674 => "001010111",
13675 => "001011110",
13676 => "001011111",
13677 => "001010111",
13678 => "001001101",
13679 => "001010110",
13680 => "001011100",
13681 => "001011100",
13682 => "001010011",
13683 => "001010010",
13684 => "001010110",
13685 => "001010111",
13686 => "001011000",
13687 => "001010011",
13688 => "001001010",
13689 => "001010110",
13690 => "001011100",
13691 => "001011110",
13692 => "001011000",
13693 => "001011100",
13694 => "001011100",
13695 => "001001111",
13696 => "001011011",
13697 => "001011011",
13698 => "001011100",
13699 => "001001110",
13700 => "001011001",
13701 => "001010110",
13702 => "001011011",
13703 => "001010000",
13704 => "001001001",
13705 => "001000110",
13706 => "001001011",
13707 => "001001000",
13708 => "000110101",
13709 => "001010001",
13710 => "001000010",
13711 => "001010110",
13712 => "001010101",
13713 => "001011001",
13714 => "001011100",
13715 => "001010101",
13716 => "001010000",
13717 => "001001110",
13718 => "001001111",
13719 => "001011001",
13720 => "001100010",
13721 => "001011010",
13722 => "001100010",
13723 => "001101101",
13724 => "001101011",
13725 => "001101111",
13726 => "001101010",
13727 => "001100001",
13728 => "001011110",
13729 => "001011000",
13730 => "001010110",
13731 => "001101010",
13732 => "000111101",
13733 => "001101101",
13734 => "001001100",
13735 => "001001111",
13736 => "001101100",
13737 => "001001000",
13738 => "001000010",
13739 => "001000110",
13740 => "000101111",
13741 => "000100100",
13742 => "000100001",
13743 => "000110111",
13744 => "001000011",
13745 => "001001010",
13746 => "000100100",
13747 => "001001001",
13748 => "001010001",
13749 => "001010011",
13750 => "001001101",
13751 => "001101011",
13752 => "001101011",
13753 => "001110010",
13754 => "001100100",
13755 => "001101100",
13756 => "001100101",
13757 => "001101110",
13758 => "001100100",
13759 => "001100001",
13760 => "001010100",
13761 => "001010000",
13762 => "001011011",
13763 => "001011001",
13764 => "001010010",
13765 => "001101101",
13766 => "001101000",
13767 => "001011100",
13768 => "001011111",
13769 => "001011100",
13770 => "001100011",
13771 => "001011000",
13772 => "001010111",
13773 => "001011100",
13774 => "001100011",
13775 => "001011011",
13776 => "001011010",
13777 => "001011100",
13778 => "001100000",
13779 => "001011011",
13780 => "001011110",
13781 => "001011110",
13782 => "001011111",
13783 => "001011001",
13784 => "001011011",
13785 => "001011111",
13786 => "001011010",
13787 => "001011000",
13788 => "001011011",
13789 => "001011000",
13790 => "001011011",
13791 => "001011110",
13792 => "001011101",
13793 => "001010011",
13794 => "001001110",
13795 => "001001111",
13796 => "001001001",
13797 => "001010010",
13798 => "001011010",
13799 => "001100011",
13800 => "001011010",
13801 => "001010111",
13802 => "001011101",
13803 => "001011011",
13804 => "001011000",
13805 => "001011110",
13806 => "001010101",
13807 => "001010000",
13808 => "001001010",
13809 => "001100011",
13810 => "001011101",
13811 => "001011111",
13812 => "001101000",
13813 => "001100100",
13814 => "001011111",
13815 => "001010110",
13816 => "001011001",
13817 => "001010111",
13818 => "001011010",
13819 => "001011000",
13820 => "001011011",
13821 => "001001110",
13822 => "001010100",
13823 => "001001111",
13824 => "001011010",
13825 => "001011001",
13826 => "001011010",
13827 => "001100000",
13828 => "001011100",
13829 => "001010100",
13830 => "001011001",
13831 => "001010110",
13832 => "001001001",
13833 => "001000110",
13834 => "001001001",
13835 => "000111111",
13836 => "001001101",
13837 => "001000001",
13838 => "001000110",
13839 => "001001100",
13840 => "001001100",
13841 => "001010101",
13842 => "001011100",
13843 => "001010010",
13844 => "001001111",
13845 => "001000000",
13846 => "000111010",
13847 => "001000000",
13848 => "001011001",
13849 => "001100010",
13850 => "001011111",
13851 => "001011100",
13852 => "001100101",
13853 => "001100011",
13854 => "001100111",
13855 => "001101001",
13856 => "001101000",
13857 => "001101011",
13858 => "001101011",
13859 => "001101101",
13860 => "001100011",
13861 => "001111111",
13862 => "001011010",
13863 => "001101111",
13864 => "001010100",
13865 => "000111111",
13866 => "001001100",
13867 => "001010101",
13868 => "001001010",
13869 => "000011110",
13870 => "000100011",
13871 => "000011110",
13872 => "000110100",
13873 => "001110001",
13874 => "001110011",
13875 => "000110010",
13876 => "000111100",
13877 => "001000010",
13878 => "001001101",
13879 => "001100011",
13880 => "001100001",
13881 => "001111000",
13882 => "001011010",
13883 => "001101111",
13884 => "001101001",
13885 => "001100010",
13886 => "001010010",
13887 => "001011010",
13888 => "001001111",
13889 => "001101100",
13890 => "001010110",
13891 => "001011000",
13892 => "001010110",
13893 => "001101111",
13894 => "001100000",
13895 => "001101000",
13896 => "001011101",
13897 => "001011101",
13898 => "001011001",
13899 => "001001101",
13900 => "001010000",
13901 => "001001110",
13902 => "001100111",
13903 => "001101100",
13904 => "001010110",
13905 => "001011111",
13906 => "001100001",
13907 => "001011100",
13908 => "001011011",
13909 => "001010111",
13910 => "001011110",
13911 => "001100101",
13912 => "001011000",
13913 => "001011100",
13914 => "001011110",
13915 => "001011100",
13916 => "001010110",
13917 => "001011100",
13918 => "001010110",
13919 => "001100010",
13920 => "001011010",
13921 => "001011110",
13922 => "001011100",
13923 => "001011011",
13924 => "001011011",
13925 => "001011001",
13926 => "001001101",
13927 => "001100011",
13928 => "001011000",
13929 => "001011001",
13930 => "001010111",
13931 => "001011101",
13932 => "001010111",
13933 => "001010110",
13934 => "001011010",
13935 => "001011000",
13936 => "001010000",
13937 => "001010001",
13938 => "001011010",
13939 => "001011010",
13940 => "001011001",
13941 => "001010101",
13942 => "001011001",
13943 => "001011011",
13944 => "001010110",
13945 => "001011000",
13946 => "001011010",
13947 => "001011100",
13948 => "001010000",
13949 => "001001111",
13950 => "001010100",
13951 => "001010010",
13952 => "001010100",
13953 => "001010011",
13954 => "001011010",
13955 => "001011101",
13956 => "001100000",
13957 => "001011000",
13958 => "001010100",
13959 => "001011110",
13960 => "001010001",
13961 => "001011110",
13962 => "001010001",
13963 => "001000001",
13964 => "001010000",
13965 => "001001001",
13966 => "000111111",
13967 => "001001001",
13968 => "001001110",
13969 => "001010101",
13970 => "001100101",
13971 => "001100010",
13972 => "001011001",
13973 => "001010001",
13974 => "001000011",
13975 => "001000000",
13976 => "001000011",
13977 => "001001111",
13978 => "001010110",
13979 => "001011110",
13980 => "001010110",
13981 => "001011110",
13982 => "001011111",
13983 => "001100000",
13984 => "001100110",
13985 => "001101001",
13986 => "001100101",
13987 => "001100111",
13988 => "001100110",
13989 => "001100111",
13990 => "001101100",
13991 => "001011101",
13992 => "001101100",
13993 => "001010100",
13994 => "001001001",
13995 => "001101010",
13996 => "001000001",
13997 => "000011010",
13998 => "000101011",
13999 => "000110100",
14000 => "001010011",
14001 => "001000101",
14002 => "001010110",
14003 => "001110011",
14004 => "000101001",
14005 => "001000011",
14006 => "001001100",
14007 => "001101110",
14008 => "010010010",
14009 => "010000110",
14010 => "001110110",
14011 => "001110100",
14012 => "001011101",
14013 => "001100111",
14014 => "001011010",
14015 => "001011101",
14016 => "001100101",
14017 => "001011110",
14018 => "001101100",
14019 => "001011001",
14020 => "001100101",
14021 => "001010110",
14022 => "001011111",
14023 => "001100101",
14024 => "001100010",
14025 => "001100001",
14026 => "001011101",
14027 => "001011010",
14028 => "001011100",
14029 => "001010111",
14030 => "001011111",
14031 => "001011110",
14032 => "001100100",
14033 => "001100010",
14034 => "001100001",
14035 => "001011010",
14036 => "001011011",
14037 => "001011000",
14038 => "001011100",
14039 => "001100101",
14040 => "001100010",
14041 => "001011101",
14042 => "001011011",
14043 => "001100000",
14044 => "001010001",
14045 => "001010101",
14046 => "001011110",
14047 => "001100101",
14048 => "001010010",
14049 => "001011100",
14050 => "001011000",
14051 => "001010001",
14052 => "001011011",
14053 => "001011011",
14054 => "001010111",
14055 => "001001010",
14056 => "001010000",
14057 => "001010001",
14058 => "001011010",
14059 => "001010001",
14060 => "001011001",
14061 => "001011000",
14062 => "001001111",
14063 => "001001110",
14064 => "001010110",
14065 => "001010111",
14066 => "001011001",
14067 => "001010110",
14068 => "001011000",
14069 => "001010010",
14070 => "001010001",
14071 => "001010011",
14072 => "001010100",
14073 => "001010110",
14074 => "001010111",
14075 => "001011001",
14076 => "001011100",
14077 => "001010101",
14078 => "001001111",
14079 => "001011000",
14080 => "001010011",
14081 => "001010100",
14082 => "001010110",
14083 => "001011010",
14084 => "001100000",
14085 => "001011100",
14086 => "001010111",
14087 => "001011101",
14088 => "001011010",
14089 => "001010000",
14090 => "001100100",
14091 => "001001101",
14092 => "001001111",
14093 => "001001110",
14094 => "001001011",
14095 => "001001111",
14096 => "001010010",
14097 => "001010000",
14098 => "001011100",
14099 => "001100001",
14100 => "001011101",
14101 => "001010101",
14102 => "001010100",
14103 => "001001001",
14104 => "000110110",
14105 => "000111011",
14106 => "000111010",
14107 => "001010111",
14108 => "001010100",
14109 => "001010100",
14110 => "001011111",
14111 => "001010101",
14112 => "001010011",
14113 => "001100101",
14114 => "001101000",
14115 => "001101000",
14116 => "001100100",
14117 => "001100011",
14118 => "001110110",
14119 => "001100000",
14120 => "001011011",
14121 => "001100111",
14122 => "001011011",
14123 => "001100110",
14124 => "001101011",
14125 => "000110000",
14126 => "001111101",
14127 => "001010010",
14128 => "000110100",
14129 => "000100010",
14130 => "000111000",
14131 => "001011101",
14132 => "001000101",
14133 => "000100111",
14134 => "000111010",
14135 => "001100011",
14136 => "001010011",
14137 => "001100001",
14138 => "001111000",
14139 => "010000000",
14140 => "010010010",
14141 => "001100100",
14142 => "001111101",
14143 => "010001010",
14144 => "001111000",
14145 => "001011111",
14146 => "001101101",
14147 => "010011011",
14148 => "001111011",
14149 => "001101100",
14150 => "001100011",
14151 => "001011101",
14152 => "001011101",
14153 => "001100110",
14154 => "001011111",
14155 => "001100001",
14156 => "001100011",
14157 => "001011010",
14158 => "001011010",
14159 => "001001011",
14160 => "001010111",
14161 => "001011111",
14162 => "001011001",
14163 => "001011010",
14164 => "001011101",
14165 => "001011111",
14166 => "001011100",
14167 => "001100011",
14168 => "001011110",
14169 => "001010000",
14170 => "001011001",
14171 => "001001101",
14172 => "001011011",
14173 => "001011000",
14174 => "001010100",
14175 => "001011011",
14176 => "001011101",
14177 => "001010110",
14178 => "001100101",
14179 => "001011000",
14180 => "001010100",
14181 => "001011001",
14182 => "001011110",
14183 => "001010110",
14184 => "001001110",
14185 => "001001001",
14186 => "001001001",
14187 => "001010011",
14188 => "001010110",
14189 => "001100101",
14190 => "001100011",
14191 => "001001110",
14192 => "000111101",
14193 => "001001110",
14194 => "001010011",
14195 => "001001111",
14196 => "001011010",
14197 => "001011100",
14198 => "001010011",
14199 => "001001111",
14200 => "001001101",
14201 => "001010001",
14202 => "001001111",
14203 => "001001010",
14204 => "001001010",
14205 => "001010011",
14206 => "001001111",
14207 => "001010001",
14208 => "001001011",
14209 => "001001100",
14210 => "001001011",
14211 => "001011010",
14212 => "001011110",
14213 => "001011001",
14214 => "001100000",
14215 => "001010111",
14216 => "001010010",
14217 => "001010101",
14218 => "001011111",
14219 => "001010001",
14220 => "001011100",
14221 => "001100000",
14222 => "001010000",
14223 => "001001100",
14224 => "001001010",
14225 => "001010111",
14226 => "001001110",
14227 => "001011110",
14228 => "001011101",
14229 => "001100000",
14230 => "001010111",
14231 => "001011000",
14232 => "001001000",
14233 => "001000011",
14234 => "000110001",
14235 => "000111100",
14236 => "001001110",
14237 => "001010100",
14238 => "001000110",
14239 => "001001110",
14240 => "000110100",
14241 => "001000010",
14242 => "001100011",
14243 => "001110011",
14244 => "001100110",
14245 => "001100111",
14246 => "001101001",
14247 => "001101001",
14248 => "001100111",
14249 => "001101100",
14250 => "001011000",
14251 => "001100110",
14252 => "001110101",
14253 => "001011101",
14254 => "001111000",
14255 => "001111010",
14256 => "001101110",
14257 => "000011001",
14258 => "000011011",
14259 => "000110111",
14260 => "001001100",
14261 => "000110011",
14262 => "001001100",
14263 => "001000110",
14264 => "001000100",
14265 => "001100010",
14266 => "001001111",
14267 => "010001011",
14268 => "010000001",
14269 => "010001010",
14270 => "001011011",
14271 => "010000011",
14272 => "001110100",
14273 => "001010100",
14274 => "001100111",
14275 => "010000001",
14276 => "001110010",
14277 => "010000100",
14278 => "001101111",
14279 => "001101000",
14280 => "001101000",
14281 => "001010001",
14282 => "001011000",
14283 => "001011001",
14284 => "001011100",
14285 => "001100000",
14286 => "001100011",
14287 => "001001111",
14288 => "001001110",
14289 => "001011110",
14290 => "001010001",
14291 => "001011001",
14292 => "001010110",
14293 => "001010001",
14294 => "001010111",
14295 => "001011100",
14296 => "001100101",
14297 => "001101100",
14298 => "001011110",
14299 => "001011110",
14300 => "001011011",
14301 => "001011101",
14302 => "001011111",
14303 => "001011001",
14304 => "001011011",
14305 => "001011001",
14306 => "001011010",
14307 => "001010101",
14308 => "001010010",
14309 => "001011010",
14310 => "001010101",
14311 => "001100001",
14312 => "001001010",
14313 => "001000111",
14314 => "001000011",
14315 => "001001000",
14316 => "001010001",
14317 => "001010111",
14318 => "001011010",
14319 => "001111000",
14320 => "001100100",
14321 => "001001100",
14322 => "001001011",
14323 => "001001010",
14324 => "001010000",
14325 => "001010100",
14326 => "001010011",
14327 => "001010100",
14328 => "001010001",
14329 => "001010010",
14330 => "001010011",
14331 => "001010010",
14332 => "001001000",
14333 => "001001001",
14334 => "001010101",
14335 => "001010100",
14336 => "001010111",
14337 => "001010100",
14338 => "001000111",
14339 => "001010111",
14340 => "001001111",
14341 => "001001110",
14342 => "001011000",
14343 => "001010011",
14344 => "001011100",
14345 => "001011100",
14346 => "001011100",
14347 => "001011100",
14348 => "001100101",
14349 => "001100011",
14350 => "001100100",
14351 => "001011001",
14352 => "001001000",
14353 => "001010011",
14354 => "001010011",
14355 => "001010101",
14356 => "001010010",
14357 => "001010011",
14358 => "001011000",
14359 => "001011101",
14360 => "001001111",
14361 => "000111110",
14362 => "001100001",
14363 => "001000000",
14364 => "000111001",
14365 => "001001111",
14366 => "001000011",
14367 => "001000001",
14368 => "001000101",
14369 => "000111001",
14370 => "001011100",
14371 => "001101010",
14372 => "001101111",
14373 => "001100010",
14374 => "001100010",
14375 => "001101010",
14376 => "001101001",
14377 => "001110000",
14378 => "001101011",
14379 => "001101101",
14380 => "001111011",
14381 => "001101010",
14382 => "001101000",
14383 => "001000010",
14384 => "000111101",
14385 => "000111001",
14386 => "000101010",
14387 => "000100001",
14388 => "001001001",
14389 => "010000101",
14390 => "001011011",
14391 => "001011100",
14392 => "001011110",
14393 => "001000001",
14394 => "001000100",
14395 => "001101110",
14396 => "001110100",
14397 => "010001010",
14398 => "001101110",
14399 => "010000100",
14400 => "001101100",
14401 => "000111110",
14402 => "000110110",
14403 => "001011011",
14404 => "000111000",
14405 => "001110111",
14406 => "001101100",
14407 => "010001100",
14408 => "010011110",
14409 => "001101110",
14410 => "001010011",
14411 => "001011010",
14412 => "001011100",
14413 => "001001011",
14414 => "001011010",
14415 => "001100000",
14416 => "001100001",
14417 => "001010110",
14418 => "001010110",
14419 => "001100110",
14420 => "001010101",
14421 => "001010100",
14422 => "001011001",
14423 => "001100000",
14424 => "001100101",
14425 => "001011111",
14426 => "001011010",
14427 => "001011101",
14428 => "001100001",
14429 => "001100001",
14430 => "001100000",
14431 => "001100000",
14432 => "001100000",
14433 => "001100100",
14434 => "001010111",
14435 => "001010000",
14436 => "001010100",
14437 => "001010110",
14438 => "001100011",
14439 => "001010101",
14440 => "001001001",
14441 => "001001010",
14442 => "001001001",
14443 => "001011001",
14444 => "001011000",
14445 => "001010110",
14446 => "001011101",
14447 => "001010101",
14448 => "001101111",
14449 => "001011111",
14450 => "001010110",
14451 => "001010111",
14452 => "001011000",
14453 => "001011110",
14454 => "001010001",
14455 => "001010001",
14456 => "001001100",
14457 => "001010101",
14458 => "001010011",
14459 => "001001001",
14460 => "001010001",
14461 => "001010011",
14462 => "001011001",
14463 => "001100101",
14464 => "001001101",
14465 => "001010001",
14466 => "001000011",
14467 => "001000101",
14468 => "001010001",
14469 => "001010001",
14470 => "001011010",
14471 => "001001110",
14472 => "001010011",
14473 => "001011101",
14474 => "001011110",
14475 => "001100000",
14476 => "001011100",
14477 => "001100010",
14478 => "001100011",
14479 => "001100000",
14480 => "001010101",
14481 => "001010001",
14482 => "001010110",
14483 => "001001011",
14484 => "001010011",
14485 => "001001100",
14486 => "001001110",
14487 => "001001000",
14488 => "001011101",
14489 => "001010001",
14490 => "001001110",
14491 => "001010100",
14492 => "001001101",
14493 => "001001000",
14494 => "001001001",
14495 => "001010000",
14496 => "001000111",
14497 => "001000010",
14498 => "001000101",
14499 => "001010100",
14500 => "001100100",
14501 => "001100000",
14502 => "001100101",
14503 => "001100111",
14504 => "001101100",
14505 => "001100100",
14506 => "001100110",
14507 => "001101101",
14508 => "001101011",
14509 => "001110011",
14510 => "001011111",
14511 => "001000011",
14512 => "001001000",
14513 => "000111111",
14514 => "000101011",
14515 => "000100100",
14516 => "000111101",
14517 => "001011001",
14518 => "001000010",
14519 => "000110010",
14520 => "001100101",
14521 => "001010110",
14522 => "001111101",
14523 => "001100111",
14524 => "001001001",
14525 => "010001101",
14526 => "010010100",
14527 => "001011000",
14528 => "001010011",
14529 => "001001001",
14530 => "000111000",
14531 => "001100111",
14532 => "001000011",
14533 => "001100001",
14534 => "001001000",
14535 => "010001011",
14536 => "010000011",
14537 => "010010010",
14538 => "001111001",
14539 => "001011010",
14540 => "001011100",
14541 => "001010101",
14542 => "001010111",
14543 => "001011001",
14544 => "001000110",
14545 => "001010110",
14546 => "001010100",
14547 => "001110000",
14548 => "001100010",
14549 => "001011111",
14550 => "001011011",
14551 => "001010101",
14552 => "001010111",
14553 => "001010101",
14554 => "001011001",
14555 => "001011011",
14556 => "001010011",
14557 => "001011100",
14558 => "001100011",
14559 => "001100001",
14560 => "001011101",
14561 => "001010101",
14562 => "001010101",
14563 => "001011000",
14564 => "001001011",
14565 => "001001010",
14566 => "001001110",
14567 => "001010110",
14568 => "001010010",
14569 => "001010101",
14570 => "001010011",
14571 => "001011001",
14572 => "001100011",
14573 => "001011010",
14574 => "001001010",
14575 => "001000001",
14576 => "001001010",
14577 => "001001111",
14578 => "001001111",
14579 => "001010000",
14580 => "001011111",
14581 => "001010001",
14582 => "001001100",
14583 => "001010100",
14584 => "001011000",
14585 => "001001001",
14586 => "001000101",
14587 => "001000001",
14588 => "001000100",
14589 => "001000101",
14590 => "001000001",
14591 => "001001010",
14592 => "001010010",
14593 => "001001010",
14594 => "001001010",
14595 => "001001110",
14596 => "001001101",
14597 => "001010011",
14598 => "001010011",
14599 => "001010100",
14600 => "001001110",
14601 => "001010111",
14602 => "001011110",
14603 => "001100010",
14604 => "001010111",
14605 => "001011101",
14606 => "001011110",
14607 => "001011111",
14608 => "001011100",
14609 => "001011010",
14610 => "001011001",
14611 => "001010111",
14612 => "001001101",
14613 => "001000110",
14614 => "001010110",
14615 => "001110001",
14616 => "001010111",
14617 => "001011100",
14618 => "001010101",
14619 => "001011010",
14620 => "001010001",
14621 => "001010000",
14622 => "001001111",
14623 => "001011101",
14624 => "001010101",
14625 => "001001011",
14626 => "001001111",
14627 => "001000110",
14628 => "001010010",
14629 => "001001101",
14630 => "001011010",
14631 => "001001110",
14632 => "001100000",
14633 => "001100101",
14634 => "001101100",
14635 => "001101100",
14636 => "001101111",
14637 => "001100100",
14638 => "001100110",
14639 => "001101101",
14640 => "001010110",
14641 => "001101000",
14642 => "000100101",
14643 => "000101111",
14644 => "000111000",
14645 => "001011111",
14646 => "001010011",
14647 => "000111001",
14648 => "001011001",
14649 => "001000100",
14650 => "001011111",
14651 => "001101011",
14652 => "001101000",
14653 => "001010000",
14654 => "001100110",
14655 => "001110001",
14656 => "001110011",
14657 => "010001101",
14658 => "001110000",
14659 => "001011001",
14660 => "001111000",
14661 => "001110100",
14662 => "010000111",
14663 => "010000001",
14664 => "001101110",
14665 => "010000000",
14666 => "010010101",
14667 => "001011010",
14668 => "001100000",
14669 => "001011100",
14670 => "000101100",
14671 => "000100010",
14672 => "001000110",
14673 => "001011111",
14674 => "001100011",
14675 => "001010000",
14676 => "001111100",
14677 => "001101100",
14678 => "001100101",
14679 => "001011100",
14680 => "001010101",
14681 => "001001110",
14682 => "001000101",
14683 => "001010000",
14684 => "001010010",
14685 => "001100111",
14686 => "001010101",
14687 => "001011011",
14688 => "001011100",
14689 => "001011011",
14690 => "001010111",
14691 => "001011111",
14692 => "001010011",
14693 => "001010010",
14694 => "001001110",
14695 => "001001011",
14696 => "001010111",
14697 => "001001110",
14698 => "001010011",
14699 => "001010101",
14700 => "001100010",
14701 => "001010100",
14702 => "001011000",
14703 => "001001110",
14704 => "001001011",
14705 => "000111111",
14706 => "001001101",
14707 => "001010001",
14708 => "001010011",
14709 => "001001010",
14710 => "001000001",
14711 => "001010011",
14712 => "001000111",
14713 => "000111111",
14714 => "001001010",
14715 => "001001010",
14716 => "001000110",
14717 => "000111111",
14718 => "001001001",
14719 => "001001111",
14720 => "001010111",
14721 => "001001111",
14722 => "001000111",
14723 => "001000011",
14724 => "001000011",
14725 => "000111111",
14726 => "001011100",
14727 => "001001011",
14728 => "001001101",
14729 => "001010000",
14730 => "001011001",
14731 => "001011000",
14732 => "001010111",
14733 => "001011111",
14734 => "001011100",
14735 => "001011101",
14736 => "001011111",
14737 => "001011010",
14738 => "001010011",
14739 => "001100100",
14740 => "001011010",
14741 => "001010000",
14742 => "001010000",
14743 => "001001100",
14744 => "001011111",
14745 => "001011101",
14746 => "001010101",
14747 => "001011011",
14748 => "001011101",
14749 => "001011001",
14750 => "001010110",
14751 => "001010111",
14752 => "001011101",
14753 => "001011111",
14754 => "001011010",
14755 => "001010001",
14756 => "001001010",
14757 => "001011101",
14758 => "001001111",
14759 => "001000100",
14760 => "001010100",
14761 => "001010011",
14762 => "001100011",
14763 => "001100100",
14764 => "001101110",
14765 => "001101011",
14766 => "001101011",
14767 => "001101001",
14768 => "001101111",
14769 => "001110001",
14770 => "001010010",
14771 => "000110101",
14772 => "000100111",
14773 => "000101011",
14774 => "000101000",
14775 => "000101010",
14776 => "001000001",
14777 => "001101000",
14778 => "001101110",
14779 => "000101111",
14780 => "001000000",
14781 => "001110110",
14782 => "001110110",
14783 => "010000001",
14784 => "010001010",
14785 => "001011010",
14786 => "001001110",
14787 => "001001101",
14788 => "000100010",
14789 => "001001110",
14790 => "001001001",
14791 => "010000011",
14792 => "010000001",
14793 => "001100001",
14794 => "001110011",
14795 => "001111101",
14796 => "001100111",
14797 => "001011000",
14798 => "001001111",
14799 => "000100011",
14800 => "000101100",
14801 => "001011000",
14802 => "001000100",
14803 => "001001001",
14804 => "001101010",
14805 => "001100010",
14806 => "001100010",
14807 => "001100000",
14808 => "001011100",
14809 => "001010001",
14810 => "001001111",
14811 => "001010111",
14812 => "001011111",
14813 => "001011100",
14814 => "001010000",
14815 => "001011101",
14816 => "001000101",
14817 => "001010011",
14818 => "001011110",
14819 => "001010010",
14820 => "001010111",
14821 => "001011000",
14822 => "001010100",
14823 => "001011011",
14824 => "001010100",
14825 => "001001110",
14826 => "001001000",
14827 => "001001011",
14828 => "001011110",
14829 => "001011111",
14830 => "001011010",
14831 => "001001111",
14832 => "001000011",
14833 => "001001001",
14834 => "001000101",
14835 => "001010101",
14836 => "001010101",
14837 => "001001100",
14838 => "001001001",
14839 => "001010011",
14840 => "001000011",
14841 => "001000101",
14842 => "001000001",
14843 => "001001010",
14844 => "001010101",
14845 => "001010001",
14846 => "001001001",
14847 => "001010000",
14848 => "001011011",
14849 => "001010111",
14850 => "001001010",
14851 => "001000010",
14852 => "001000011",
14853 => "001001101",
14854 => "001100110",
14855 => "001010011",
14856 => "001001101",
14857 => "001010101",
14858 => "001011111",
14859 => "001011000",
14860 => "001100110",
14861 => "001101010",
14862 => "001100010",
14863 => "001010001",
14864 => "001010101",
14865 => "001100001",
14866 => "001101000",
14867 => "001011000",
14868 => "001010100",
14869 => "001010011",
14870 => "001010011",
14871 => "001010100",
14872 => "001011110",
14873 => "001010111",
14874 => "001010110",
14875 => "001101110",
14876 => "001101001",
14877 => "001010110",
14878 => "001011100",
14879 => "001011011",
14880 => "001011101",
14881 => "001100001",
14882 => "001100100",
14883 => "001011010",
14884 => "001100001",
14885 => "001101000",
14886 => "001011001",
14887 => "001011000",
14888 => "001011101",
14889 => "001100011",
14890 => "001100100",
14891 => "001011101",
14892 => "001101000",
14893 => "001100001",
14894 => "001010111",
14895 => "001100000",
14896 => "001011110",
14897 => "001101111",
14898 => "001100100",
14899 => "001010001",
14900 => "001010010",
14901 => "001001111",
14902 => "000110110",
14903 => "000100100",
14904 => "001000001",
14905 => "001000110",
14906 => "001000100",
14907 => "001100110",
14908 => "000101101",
14909 => "010000000",
14910 => "001100001",
14911 => "001110011",
14912 => "001101011",
14913 => "001011100",
14914 => "000111101",
14915 => "000101101",
14916 => "000011011",
14917 => "000101111",
14918 => "001010001",
14919 => "000111001",
14920 => "000101111",
14921 => "001100010",
14922 => "001101101",
14923 => "001101010",
14924 => "001100001",
14925 => "001000110",
14926 => "001100101",
14927 => "001001001",
14928 => "000110111",
14929 => "000100011",
14930 => "001000001",
14931 => "001000001",
14932 => "001010110",
14933 => "001100101",
14934 => "001100000",
14935 => "001100001",
14936 => "001100010",
14937 => "001010011",
14938 => "001001110",
14939 => "001001101",
14940 => "001010110",
14941 => "001010101",
14942 => "001100000",
14943 => "001011110",
14944 => "001011000",
14945 => "001010011",
14946 => "001011001",
14947 => "001011010",
14948 => "001011101",
14949 => "001011100",
14950 => "001100010",
14951 => "001011101",
14952 => "001010101",
14953 => "001010001",
14954 => "001001111",
14955 => "001001110",
14956 => "001010110",
14957 => "001011110",
14958 => "001010100",
14959 => "001010100",
14960 => "001010011",
14961 => "001000110",
14962 => "001000011",
14963 => "001001110",
14964 => "001010011",
14965 => "001001011",
14966 => "001001110",
14967 => "001000110",
14968 => "001000000",
14969 => "001000010",
14970 => "001001011",
14971 => "001001010",
14972 => "001011100",
14973 => "001001010",
14974 => "001001001",
14975 => "001010010",
14976 => "001010110",
14977 => "001010101",
14978 => "001001011",
14979 => "001001111",
14980 => "001010110",
14981 => "001001100",
14982 => "001001111",
14983 => "001000111",
14984 => "001010011",
14985 => "001010010",
14986 => "001010010",
14987 => "001100010",
14988 => "001100001",
14989 => "001011110",
14990 => "001011100",
14991 => "001011010",
14992 => "001010111",
14993 => "001100001",
14994 => "001011110",
14995 => "001100100",
14996 => "001100000",
14997 => "001011100",
14998 => "001011000",
14999 => "001001101",
15000 => "001010000",
15001 => "001010101",
15002 => "001011000",
15003 => "001011110",
15004 => "001100111",
15005 => "001010110",
15006 => "001010001",
15007 => "001011010",
15008 => "001011110",
15009 => "001011001",
15010 => "001100101",
15011 => "001011100",
15012 => "001100101",
15013 => "001010011",
15014 => "001011001",
15015 => "001100000",
15016 => "001100100",
15017 => "001100010",
15018 => "001100101",
15019 => "001101110",
15020 => "001100010",
15021 => "001011011",
15022 => "001000111",
15023 => "001001010",
15024 => "001010110",
15025 => "001101000",
15026 => "001110100",
15027 => "001101001",
15028 => "001000111",
15029 => "001001110",
15030 => "000101001",
15031 => "000100000",
15032 => "000110111",
15033 => "000110010",
15034 => "001101101",
15035 => "001101000",
15036 => "001001101",
15037 => "001010001",
15038 => "001111101",
15039 => "010010101",
15040 => "000111000",
15041 => "001010011",
15042 => "001101111",
15043 => "000010011",
15044 => "000011010",
15045 => "000101100",
15046 => "000101011",
15047 => "000110101",
15048 => "001010111",
15049 => "001101011",
15050 => "001111010",
15051 => "001011110",
15052 => "001000010",
15053 => "001000110",
15054 => "001001010",
15055 => "001001010",
15056 => "000110010",
15057 => "000101011",
15058 => "001010010",
15059 => "000110000",
15060 => "001000110",
15061 => "001011110",
15062 => "001100010",
15063 => "001011011",
15064 => "001100011",
15065 => "001100011",
15066 => "001011111",
15067 => "001011011",
15068 => "001100000",
15069 => "001011010",
15070 => "001011010",
15071 => "001010101",
15072 => "001010111",
15073 => "001011010",
15074 => "001010110",
15075 => "001011101",
15076 => "001001101",
15077 => "001100100",
15078 => "001101101",
15079 => "001100110",
15080 => "001011110",
15081 => "001010001",
15082 => "001010001",
15083 => "001001001",
15084 => "001001100",
15085 => "001001110",
15086 => "001010101",
15087 => "001001101",
15088 => "001000110",
15089 => "001010001",
15090 => "001001010",
15091 => "001000110",
15092 => "001000010",
15093 => "001010000",
15094 => "001001110",
15095 => "001010001",
15096 => "001011110",
15097 => "001001000",
15098 => "001000101",
15099 => "001000101",
15100 => "001001001",
15101 => "001001010",
15102 => "001000010",
15103 => "000110101",
15104 => "001010010",
15105 => "001001111",
15106 => "001001110",
15107 => "001011010",
15108 => "001010000",
15109 => "001010011",
15110 => "001001101",
15111 => "001001101",
15112 => "001001010",
15113 => "001000110",
15114 => "001011010",
15115 => "001100110",
15116 => "001011111",
15117 => "001011010",
15118 => "001011000",
15119 => "001011001",
15120 => "001010011",
15121 => "001010000",
15122 => "001010111",
15123 => "001011101",
15124 => "001011111",
15125 => "001100011",
15126 => "001011111",
15127 => "001011110",
15128 => "001100100",
15129 => "001100000",
15130 => "001010111",
15131 => "001100010",
15132 => "001010010",
15133 => "001010011",
15134 => "001001011",
15135 => "001010110",
15136 => "001010111",
15137 => "001011000",
15138 => "001100010",
15139 => "001101101",
15140 => "001011110",
15141 => "001010110",
15142 => "001001100",
15143 => "001010100",
15144 => "001011111",
15145 => "001011111",
15146 => "001011011",
15147 => "001100011",
15148 => "001011011",
15149 => "001010110",
15150 => "001010110",
15151 => "001010010",
15152 => "001011001",
15153 => "001010111",
15154 => "001100111",
15155 => "001101000",
15156 => "001101101",
15157 => "001011000",
15158 => "001001011",
15159 => "000110111",
15160 => "001010110",
15161 => "000111000",
15162 => "000110010",
15163 => "001001001",
15164 => "001100100",
15165 => "001000010",
15166 => "001001101",
15167 => "000110101",
15168 => "001100111",
15169 => "000111011",
15170 => "000111011",
15171 => "000111100",
15172 => "000001011",
15173 => "000111101",
15174 => "000010111",
15175 => "000101000",
15176 => "000110000",
15177 => "000111100",
15178 => "001010110",
15179 => "001010111",
15180 => "001011100",
15181 => "001101001",
15182 => "000110101",
15183 => "000111011",
15184 => "001000001",
15185 => "000111011",
15186 => "000110101",
15187 => "000010111",
15188 => "000101100",
15189 => "001000011",
15190 => "001001100",
15191 => "001100000",
15192 => "001100000",
15193 => "001100101",
15194 => "001011010",
15195 => "001011010",
15196 => "001010101",
15197 => "001011001",
15198 => "001011000",
15199 => "001011001",
15200 => "001011100",
15201 => "001011010",
15202 => "001100010",
15203 => "001011110",
15204 => "001011101",
15205 => "001011001",
15206 => "001100000",
15207 => "001010100",
15208 => "001011101",
15209 => "001100000",
15210 => "001011101",
15211 => "001010100",
15212 => "001001010",
15213 => "001001100",
15214 => "001001100",
15215 => "001011000",
15216 => "001100000",
15217 => "001101000",
15218 => "001010001",
15219 => "001001110",
15220 => "001001101",
15221 => "001001011",
15222 => "001001001",
15223 => "001000110",
15224 => "001001000",
15225 => "001010010",
15226 => "001001111",
15227 => "001001110",
15228 => "001000110",
15229 => "001001000",
15230 => "001001000",
15231 => "001000010",
15232 => "001001100",
15233 => "001000111",
15234 => "001001111",
15235 => "001001111",
15236 => "001001110",
15237 => "001011100",
15238 => "001011001",
15239 => "001010101",
15240 => "001001100",
15241 => "001000111",
15242 => "001001111",
15243 => "001100100",
15244 => "001011101",
15245 => "001010111",
15246 => "001011100",
15247 => "001011101",
15248 => "001010011",
15249 => "001010011",
15250 => "001001101",
15251 => "001010001",
15252 => "001011000",
15253 => "001011101",
15254 => "001011110",
15255 => "001100000",
15256 => "001100011",
15257 => "001101000",
15258 => "001100011",
15259 => "001011110",
15260 => "001010110",
15261 => "001010111",
15262 => "001001111",
15263 => "001010011",
15264 => "001010001",
15265 => "001011101",
15266 => "001100010",
15267 => "001100010",
15268 => "001011101",
15269 => "001010000",
15270 => "001000100",
15271 => "001011010",
15272 => "001011000",
15273 => "001011011",
15274 => "001010011",
15275 => "001011101",
15276 => "001011011",
15277 => "001100101",
15278 => "001100110",
15279 => "001100101",
15280 => "001011001",
15281 => "001011001",
15282 => "001100010",
15283 => "001100100",
15284 => "001100000",
15285 => "001100101",
15286 => "001101001",
15287 => "001010001",
15288 => "001010100",
15289 => "000110101",
15290 => "000110000",
15291 => "000111110",
15292 => "001001101",
15293 => "000101010",
15294 => "000101000",
15295 => "000100110",
15296 => "001001110",
15297 => "000110011",
15298 => "000011110",
15299 => "000001101",
15300 => "000001011",
15301 => "000101000",
15302 => "000100100",
15303 => "000100010",
15304 => "000100011",
15305 => "000100100",
15306 => "000101011",
15307 => "001011001",
15308 => "001001011",
15309 => "000110111",
15310 => "001010101",
15311 => "001001111",
15312 => "001000101",
15313 => "001000000",
15314 => "000110110",
15315 => "001001110",
15316 => "001001001",
15317 => "000111000",
15318 => "000111001",
15319 => "001000100",
15320 => "001001011",
15321 => "001000101",
15322 => "001100110",
15323 => "001010110",
15324 => "001001001",
15325 => "001010101",
15326 => "001010101",
15327 => "001011010",
15328 => "001010000",
15329 => "001010011",
15330 => "001010111",
15331 => "001100000",
15332 => "001100010",
15333 => "001011110",
15334 => "001001011",
15335 => "001010011",
15336 => "001011000",
15337 => "001011010",
15338 => "001010111",
15339 => "001010101",
15340 => "001010111",
15341 => "001001111",
15342 => "001010000",
15343 => "001000111",
15344 => "001001010",
15345 => "001011110",
15346 => "001101001",
15347 => "001011010",
15348 => "001011000",
15349 => "001010110",
15350 => "001010001",
15351 => "001001010",
15352 => "001001100",
15353 => "001001000",
15354 => "001000011",
15355 => "001001000",
15356 => "001001000",
15357 => "001001010",
15358 => "001010001",
15359 => "001000001",
15360 => "001010000",
15361 => "001000000",
15362 => "001001010",
15363 => "001001111",
15364 => "001101001",
15365 => "001001110",
15366 => "001010101",
15367 => "001010111",
15368 => "001011101",
15369 => "001010111",
15370 => "001001111",
15371 => "001010100",
15372 => "001011011",
15373 => "001010001",
15374 => "001001111",
15375 => "001011100",
15376 => "001011011",
15377 => "001011011",
15378 => "001011111",
15379 => "001011001",
15380 => "001011001",
15381 => "001011010",
15382 => "001010101",
15383 => "001011101",
15384 => "001100011",
15385 => "001100110",
15386 => "001011011",
15387 => "001011010",
15388 => "001011110",
15389 => "001100101",
15390 => "001011101",
15391 => "001001101",
15392 => "001011100",
15393 => "001011001",
15394 => "001001101",
15395 => "001010100",
15396 => "001010111",
15397 => "001001110",
15398 => "000111100",
15399 => "001001001",
15400 => "001010111",
15401 => "001001100",
15402 => "001010011",
15403 => "001010010",
15404 => "001010100",
15405 => "001101000",
15406 => "001011101",
15407 => "001110000",
15408 => "001100011",
15409 => "001100000",
15410 => "001100001",
15411 => "001101000",
15412 => "001011101",
15413 => "001011011",
15414 => "001101010",
15415 => "001101001",
15416 => "001100101",
15417 => "001001110",
15418 => "001000110",
15419 => "000110100",
15420 => "001000111",
15421 => "000101001",
15422 => "000010011",
15423 => "000101101",
15424 => "000100111",
15425 => "001000101",
15426 => "000111000",
15427 => "000010010",
15428 => "000001100",
15429 => "000011010",
15430 => "000001111",
15431 => "000010011",
15432 => "000001011",
15433 => "000001111",
15434 => "000100001",
15435 => "000110100",
15436 => "000100001",
15437 => "001000000",
15438 => "001010100",
15439 => "001001011",
15440 => "000101111",
15441 => "001110001",
15442 => "010001101",
15443 => "001110000",
15444 => "001001110",
15445 => "001001100",
15446 => "000111001",
15447 => "001000010",
15448 => "001001111",
15449 => "001000010",
15450 => "001001111",
15451 => "001100000",
15452 => "001100101",
15453 => "001001011",
15454 => "001011010",
15455 => "001011011",
15456 => "000111001",
15457 => "001010001",
15458 => "001001011",
15459 => "001000111",
15460 => "001100001",
15461 => "001011100",
15462 => "001010111",
15463 => "001010100",
15464 => "001011100",
15465 => "001011001",
15466 => "001011000",
15467 => "001011101",
15468 => "001011110",
15469 => "001011100",
15470 => "001011001",
15471 => "001011010",
15472 => "001010100",
15473 => "001010001",
15474 => "001010010",
15475 => "001000100",
15476 => "000111110",
15477 => "001000100",
15478 => "001001000",
15479 => "001001100",
15480 => "001010010",
15481 => "001001101",
15482 => "001010001",
15483 => "001010110",
15484 => "001001001",
15485 => "001010011",
15486 => "001010101",
15487 => "001010100",
15488 => "001001101",
15489 => "001001101",
15490 => "001001100",
15491 => "001010101",
15492 => "001100011",
15493 => "001001110",
15494 => "001011011",
15495 => "001010000",
15496 => "001011000",
15497 => "001010000",
15498 => "001010001",
15499 => "001011010",
15500 => "001011010",
15501 => "001010010",
15502 => "001100011",
15503 => "001010111",
15504 => "001010110",
15505 => "001011000",
15506 => "001011111",
15507 => "001100111",
15508 => "001001110",
15509 => "001001110",
15510 => "001001010",
15511 => "001011111",
15512 => "001011011",
15513 => "001011010",
15514 => "001010110",
15515 => "001011100",
15516 => "001011000",
15517 => "001101000",
15518 => "001010100",
15519 => "001010101",
15520 => "001010001",
15521 => "001001011",
15522 => "001001100",
15523 => "001010001",
15524 => "001010111",
15525 => "001010001",
15526 => "001001110",
15527 => "001010011",
15528 => "001001011",
15529 => "001010000",
15530 => "001001111",
15531 => "001010000",
15532 => "001011110",
15533 => "001100011",
15534 => "001100100",
15535 => "001101000",
15536 => "001101010",
15537 => "001100101",
15538 => "001100000",
15539 => "001010111",
15540 => "001010111",
15541 => "001011010",
15542 => "001011001",
15543 => "001101101",
15544 => "001011111",
15545 => "001100110",
15546 => "001010000",
15547 => "001001100",
15548 => "001010000",
15549 => "000111010",
15550 => "000111101",
15551 => "000110100",
15552 => "000110001",
15553 => "000110110",
15554 => "001000010",
15555 => "000011011",
15556 => "000010101",
15557 => "000111010",
15558 => "000100110",
15559 => "000011100",
15560 => "000001101",
15561 => "000010000",
15562 => "000010110",
15563 => "000010010",
15564 => "000110001",
15565 => "000011101",
15566 => "000110010",
15567 => "000111001",
15568 => "000110100",
15569 => "000111100",
15570 => "000101101",
15571 => "001001100",
15572 => "001001101",
15573 => "000110011",
15574 => "000111011",
15575 => "000101100",
15576 => "000111101",
15577 => "001000101",
15578 => "001000011",
15579 => "000111111",
15580 => "001010010",
15581 => "001101110",
15582 => "001100000",
15583 => "001110101",
15584 => "001011000",
15585 => "001010110",
15586 => "001010001",
15587 => "001000001",
15588 => "001011001",
15589 => "001001101",
15590 => "001010001",
15591 => "001010001",
15592 => "001010110",
15593 => "001011111",
15594 => "001011010",
15595 => "001001111",
15596 => "001011110",
15597 => "001011010",
15598 => "001011001",
15599 => "001010111",
15600 => "001100001",
15601 => "001001011",
15602 => "001001110",
15603 => "001010110",
15604 => "001001101",
15605 => "001001001",
15606 => "001001101",
15607 => "001001011",
15608 => "001010000",
15609 => "001001110",
15610 => "001010100",
15611 => "001010000",
15612 => "001010100",
15613 => "001000110",
15614 => "001001011",
15615 => "001010111",
15616 => "001000011",
15617 => "001000100",
15618 => "001000011",
15619 => "001000101",
15620 => "001011010",
15621 => "001001011",
15622 => "001001110",
15623 => "001001100",
15624 => "001010010",
15625 => "001010100",
15626 => "001010000",
15627 => "001001110",
15628 => "001010001",
15629 => "001010001",
15630 => "001011011",
15631 => "001010100",
15632 => "001011000",
15633 => "001010100",
15634 => "001011001",
15635 => "001010000",
15636 => "001001001",
15637 => "001010010",
15638 => "001001000",
15639 => "001010101",
15640 => "001011110",
15641 => "001001101",
15642 => "001011011",
15643 => "001000101",
15644 => "001001101",
15645 => "001001110",
15646 => "001001110",
15647 => "001001011",
15648 => "001011000",
15649 => "001001100",
15650 => "001011000",
15651 => "001000111",
15652 => "001001010",
15653 => "001000000",
15654 => "000111000",
15655 => "000110101",
15656 => "000111010",
15657 => "001001111",
15658 => "001001000",
15659 => "001001000",
15660 => "001010110",
15661 => "001001111",
15662 => "001100001",
15663 => "001011010",
15664 => "001101010",
15665 => "001011111",
15666 => "001011100",
15667 => "001010010",
15668 => "001010100",
15669 => "001010011",
15670 => "001001010",
15671 => "001010111",
15672 => "001011011",
15673 => "001011000",
15674 => "001101001",
15675 => "001100100",
15676 => "001101011",
15677 => "001101010",
15678 => "001011001",
15679 => "001010001",
15680 => "000111011",
15681 => "001001100",
15682 => "000101101",
15683 => "000011001",
15684 => "000000100",
15685 => "000111010",
15686 => "000101000",
15687 => "000111011",
15688 => "000001110",
15689 => "000001100",
15690 => "000100010",
15691 => "000100000",
15692 => "000100111",
15693 => "000100110",
15694 => "000110110",
15695 => "000101111",
15696 => "000011100",
15697 => "000011001",
15698 => "000011111",
15699 => "000100000",
15700 => "000100011",
15701 => "000100010",
15702 => "000100001",
15703 => "000110001",
15704 => "001000110",
15705 => "001000110",
15706 => "000111110",
15707 => "001000010",
15708 => "001001011",
15709 => "000111101",
15710 => "001000100",
15711 => "001010101",
15712 => "001100011",
15713 => "001000111",
15714 => "001001110",
15715 => "001011010",
15716 => "001101101",
15717 => "001100011",
15718 => "001010011",
15719 => "001011100",
15720 => "001011010",
15721 => "001010111",
15722 => "001010110",
15723 => "001010010",
15724 => "001011110",
15725 => "001100000",
15726 => "001011010",
15727 => "001011100",
15728 => "001011100",
15729 => "001010101",
15730 => "001001101",
15731 => "001000000",
15732 => "001000100",
15733 => "001001011",
15734 => "001010000",
15735 => "001001111",
15736 => "001001001",
15737 => "001001010",
15738 => "001010011",
15739 => "001010010",
15740 => "001010111",
15741 => "001011101",
15742 => "001010011",
15743 => "001010010",
15744 => "001000100",
15745 => "001001111",
15746 => "001000101",
15747 => "001010001",
15748 => "001001011",
15749 => "001000111",
15750 => "000111101",
15751 => "001000110",
15752 => "001010110",
15753 => "001000110",
15754 => "001000111",
15755 => "001010111",
15756 => "001011101",
15757 => "001001101",
15758 => "001010000",
15759 => "001010000",
15760 => "001010001",
15761 => "001011110",
15762 => "001100001",
15763 => "001001001",
15764 => "001000011",
15765 => "001011001",
15766 => "001010100",
15767 => "001011110",
15768 => "001011011",
15769 => "001010101",
15770 => "001010010",
15771 => "000111011",
15772 => "000110110",
15773 => "001010110",
15774 => "001000100",
15775 => "001001010",
15776 => "001001010",
15777 => "001010011",
15778 => "001000001",
15779 => "001001011",
15780 => "001010100",
15781 => "001001000",
15782 => "001000110",
15783 => "000111110",
15784 => "000110110",
15785 => "001000110",
15786 => "001000100",
15787 => "001010011",
15788 => "001010011",
15789 => "001000010",
15790 => "001010100",
15791 => "001001010",
15792 => "001011100",
15793 => "001101001",
15794 => "001100100",
15795 => "001011000",
15796 => "001001101",
15797 => "001010100",
15798 => "001001111",
15799 => "001010011",
15800 => "001010011",
15801 => "001010100",
15802 => "001100001",
15803 => "001100101",
15804 => "001101101",
15805 => "001101011",
15806 => "001011110",
15807 => "001011010",
15808 => "000100111",
15809 => "000100101",
15810 => "000010010",
15811 => "000010101",
15812 => "000010100",
15813 => "000011110",
15814 => "000111000",
15815 => "000111111",
15816 => "000100100",
15817 => "000100001",
15818 => "000010011",
15819 => "000100011",
15820 => "000010101",
15821 => "000011100",
15822 => "000011011",
15823 => "000011111",
15824 => "000011100",
15825 => "000101111",
15826 => "000101000",
15827 => "000110001",
15828 => "000100010",
15829 => "000101101",
15830 => "000010001",
15831 => "000100100",
15832 => "000110011",
15833 => "001010110",
15834 => "000111101",
15835 => "000100000",
15836 => "001000011",
15837 => "000111001",
15838 => "001000001",
15839 => "001000001",
15840 => "001001001",
15841 => "001100011",
15842 => "001000010",
15843 => "001100011",
15844 => "001011110",
15845 => "001010001",
15846 => "000111101",
15847 => "001011010",
15848 => "001100000",
15849 => "001100010",
15850 => "001011101",
15851 => "001100011",
15852 => "001011111",
15853 => "001011101",
15854 => "001011000",
15855 => "001000101",
15856 => "001000110",
15857 => "001000100",
15858 => "001010001",
15859 => "001001100",
15860 => "001000011",
15861 => "001000101",
15862 => "001011000",
15863 => "001000101",
15864 => "001010011",
15865 => "001001001",
15866 => "001000101",
15867 => "001011001",
15868 => "001000000",
15869 => "001001001",
15870 => "001001010",
15871 => "001001000",
15872 => "001000101",
15873 => "001001101",
15874 => "001001010",
15875 => "001001001",
15876 => "001001001",
15877 => "001001110",
15878 => "001001110",
15879 => "001011001",
15880 => "001001000",
15881 => "001000101",
15882 => "001000100",
15883 => "001010001",
15884 => "001011011",
15885 => "001011000",
15886 => "001001110",
15887 => "001011001",
15888 => "001010011",
15889 => "001010100",
15890 => "001011010",
15891 => "001001011",
15892 => "001001100",
15893 => "001010110",
15894 => "001001111",
15895 => "001010110",
15896 => "001010010",
15897 => "001010110",
15898 => "001000100",
15899 => "001001111",
15900 => "001011110",
15901 => "001010010",
15902 => "001001001",
15903 => "001000011",
15904 => "000111010",
15905 => "001001000",
15906 => "001001010",
15907 => "001010101",
15908 => "001001100",
15909 => "001000011",
15910 => "000111110",
15911 => "001000011",
15912 => "001000110",
15913 => "001000101",
15914 => "000111101",
15915 => "001000001",
15916 => "000111010",
15917 => "001000110",
15918 => "000111010",
15919 => "001000000",
15920 => "001010110",
15921 => "001011100",
15922 => "001011001",
15923 => "001100000",
15924 => "001011001",
15925 => "001010101",
15926 => "001001001",
15927 => "001001011",
15928 => "001001001",
15929 => "001010110",
15930 => "001100000",
15931 => "001100011",
15932 => "001011100",
15933 => "001101101",
15934 => "001100011",
15935 => "001100011",
15936 => "001010100",
15937 => "000101010",
15938 => "000011011",
15939 => "000010001",
15940 => "000010000",
15941 => "000101001",
15942 => "000111011",
15943 => "001010111",
15944 => "001001110",
15945 => "000110000",
15946 => "000110000",
15947 => "000101010",
15948 => "000011110",
15949 => "000010101",
15950 => "000100011",
15951 => "000010101",
15952 => "000010101",
15953 => "000100100",
15954 => "000101011",
15955 => "000100011",
15956 => "000011101",
15957 => "000011000",
15958 => "000001110",
15959 => "000010101",
15960 => "000010011",
15961 => "001001100",
15962 => "000100110",
15963 => "000110000",
15964 => "000110010",
15965 => "000110001",
15966 => "001011111",
15967 => "001000000",
15968 => "000110111",
15969 => "001001110",
15970 => "001001100",
15971 => "000110001",
15972 => "001011110",
15973 => "000111110",
15974 => "001010000",
15975 => "001100110",
15976 => "001100010",
15977 => "001100010",
15978 => "001011101",
15979 => "001011100",
15980 => "001011101",
15981 => "001011001",
15982 => "001011111",
15983 => "001011101",
15984 => "001010011",
15985 => "001001100",
15986 => "001010010",
15987 => "001010010",
15988 => "001001101",
15989 => "001001100",
15990 => "001001010",
15991 => "001010110",
15992 => "001010100",
15993 => "001001111",
15994 => "001001101",
15995 => "001010101",
15996 => "001000111",
15997 => "001010010",
15998 => "001010000",
15999 => "001011001",
16000 => "001000011",
16001 => "001011000",
16002 => "000111010",
16003 => "001001101",
16004 => "001001101",
16005 => "001000001",
16006 => "001000010",
16007 => "001010010",
16008 => "001001001",
16009 => "001000111",
16010 => "001010110",
16011 => "001001110",
16012 => "001001011",
16013 => "001011000",
16014 => "001100000",
16015 => "001010000",
16016 => "001011011",
16017 => "001010111",
16018 => "001001011",
16019 => "001001000",
16020 => "001001110",
16021 => "001001001",
16022 => "001010001",
16023 => "001010010",
16024 => "001001011",
16025 => "001010011",
16026 => "000111101",
16027 => "001010011",
16028 => "001010011",
16029 => "001010111",
16030 => "000111101",
16031 => "001010010",
16032 => "001001001",
16033 => "001011000",
16034 => "001011000",
16035 => "001010001",
16036 => "001000011",
16037 => "001000000",
16038 => "001000101",
16039 => "001000001",
16040 => "001001001",
16041 => "001001100",
16042 => "001001000",
16043 => "001000100",
16044 => "001000100",
16045 => "000111110",
16046 => "001000100",
16047 => "000111101",
16048 => "001001100",
16049 => "001010001",
16050 => "001011110",
16051 => "001010110",
16052 => "001010001",
16053 => "001001001",
16054 => "001001001",
16055 => "001001100",
16056 => "001010100",
16057 => "001011010",
16058 => "001011000",
16059 => "001011100",
16060 => "001010110",
16061 => "001011111",
16062 => "001101010",
16063 => "001101101",
16064 => "001101001",
16065 => "001010111",
16066 => "000110010",
16067 => "000111011",
16068 => "000100111",
16069 => "001001001",
16070 => "000101100",
16071 => "000110100",
16072 => "001001000",
16073 => "000111011",
16074 => "000111001",
16075 => "000111011",
16076 => "000110011",
16077 => "000010101",
16078 => "000011010",
16079 => "000010011",
16080 => "000010011",
16081 => "000010110",
16082 => "000110111",
16083 => "000110010",
16084 => "000101111",
16085 => "000101010",
16086 => "000010111",
16087 => "000011011",
16088 => "000001111",
16089 => "000100100",
16090 => "000100101",
16091 => "000010111",
16092 => "000101000",
16093 => "000100010",
16094 => "000110001",
16095 => "000101010",
16096 => "000110101",
16097 => "000111010",
16098 => "001000011",
16099 => "000100110",
16100 => "000110111",
16101 => "000111010",
16102 => "001100100",
16103 => "001001011",
16104 => "001011101",
16105 => "001010001",
16106 => "001011011",
16107 => "001011001",
16108 => "001100110",
16109 => "001100011",
16110 => "001011011",
16111 => "001001100",
16112 => "001001101",
16113 => "001010010",
16114 => "001010101",
16115 => "001010010",
16116 => "001001110",
16117 => "001000111",
16118 => "000111111",
16119 => "000111110",
16120 => "001000101",
16121 => "001001010",
16122 => "001001100",
16123 => "001001100",
16124 => "001001000",
16125 => "001010001",
16126 => "001000010",
16127 => "001000000",
16128 => "001001101",
16129 => "001000101",
16130 => "001001011",
16131 => "001001000",
16132 => "001000100",
16133 => "001001001",
16134 => "001010011",
16135 => "001001011",
16136 => "001001101",
16137 => "001000100",
16138 => "001001111",
16139 => "001010010",
16140 => "001001101",
16141 => "001011000",
16142 => "001011100",
16143 => "001100011",
16144 => "001011011",
16145 => "001010100",
16146 => "001010011",
16147 => "001000111",
16148 => "001010001",
16149 => "001001100",
16150 => "001010011",
16151 => "001001000",
16152 => "001011010",
16153 => "001011000",
16154 => "001010000",
16155 => "001010000",
16156 => "001010000",
16157 => "001001010",
16158 => "001000011",
16159 => "001000110",
16160 => "001001000",
16161 => "001001111",
16162 => "001010011",
16163 => "001011110",
16164 => "001011010",
16165 => "000111111",
16166 => "001001101",
16167 => "001001101",
16168 => "001001001",
16169 => "001001101",
16170 => "001010001",
16171 => "001010001",
16172 => "000111101",
16173 => "001001000",
16174 => "001000100",
16175 => "001000101",
16176 => "001001000",
16177 => "001001011",
16178 => "001000010",
16179 => "001001011",
16180 => "001010001",
16181 => "001010000",
16182 => "001010010",
16183 => "001011010",
16184 => "001011001",
16185 => "001011011",
16186 => "001011000",
16187 => "001011110",
16188 => "001100000",
16189 => "001010010",
16190 => "001010010",
16191 => "001101010",
16192 => "001111001",
16193 => "001100100",
16194 => "001100101",
16195 => "001001000",
16196 => "000111000",
16197 => "000101000",
16198 => "000011010",
16199 => "000101110",
16200 => "000011001",
16201 => "000011001",
16202 => "000100110",
16203 => "000110001",
16204 => "000100110",
16205 => "000100101",
16206 => "000101101",
16207 => "000011111",
16208 => "000011110",
16209 => "000011111",
16210 => "000100101",
16211 => "000111010",
16212 => "000111101",
16213 => "000011111",
16214 => "000110010",
16215 => "000011001",
16216 => "000010001",
16217 => "000100001",
16218 => "000101010",
16219 => "000011101",
16220 => "000110110",
16221 => "000101001",
16222 => "000101111",
16223 => "000101110",
16224 => "000101100",
16225 => "000101100",
16226 => "001001000",
16227 => "000101000",
16228 => "000111010",
16229 => "001000111",
16230 => "001011000",
16231 => "001011110",
16232 => "001101101",
16233 => "001111011",
16234 => "001011000",
16235 => "001011000",
16236 => "001011000",
16237 => "001010010",
16238 => "001011110",
16239 => "001011110",
16240 => "001001110",
16241 => "001011010",
16242 => "001011010",
16243 => "001010100",
16244 => "001010101",
16245 => "001011010",
16246 => "001010101",
16247 => "001010010",
16248 => "001001000",
16249 => "001001001",
16250 => "001001001",
16251 => "001000110",
16252 => "001000110",
16253 => "001010110",
16254 => "001011111",
16255 => "001010010",
16256 => "001001111",
16257 => "001000110",
16258 => "001000101",
16259 => "001000010",
16260 => "001001111",
16261 => "001010011",
16262 => "001001111",
16263 => "001010001",
16264 => "001001110",
16265 => "001001111",
16266 => "001000100",
16267 => "001010110",
16268 => "001001001",
16269 => "001001100",
16270 => "001010101",
16271 => "001011001",
16272 => "001011011",
16273 => "001010100",
16274 => "001010011",
16275 => "001001011",
16276 => "001011111",
16277 => "001000101",
16278 => "001001111",
16279 => "001010000",
16280 => "001010001",
16281 => "001010101",
16282 => "001001111",
16283 => "001011110",
16284 => "001001100",
16285 => "001010101",
16286 => "001010010",
16287 => "000111110",
16288 => "001000100",
16289 => "001001000",
16290 => "001001011",
16291 => "001010010",
16292 => "001011001",
16293 => "001010000",
16294 => "001010111",
16295 => "001010010",
16296 => "001100000",
16297 => "001100001",
16298 => "001011000",
16299 => "001001110",
16300 => "001010110",
16301 => "001000101",
16302 => "001000000",
16303 => "000111110",
16304 => "001001010",
16305 => "001001000",
16306 => "001001101",
16307 => "001000001",
16308 => "001010011",
16309 => "001010110",
16310 => "001011010",
16311 => "001010101",
16312 => "001010101",
16313 => "001011000",
16314 => "001010100",
16315 => "001010101",
16316 => "001010110",
16317 => "001011101",
16318 => "001011100",
16319 => "001011010",
16320 => "001010011",
16321 => "001100110",
16322 => "001100010",
16323 => "001011101",
16324 => "001011000",
16325 => "001001010",
16326 => "001010001",
16327 => "001000000",
16328 => "000100101",
16329 => "000100101",
16330 => "000101100",
16331 => "000110011",
16332 => "000101010",
16333 => "000101001",
16334 => "000100110",
16335 => "000100011",
16336 => "000100010",
16337 => "000111011",
16338 => "000101010",
16339 => "000110111",
16340 => "001001100",
16341 => "000111110",
16342 => "000111010",
16343 => "000101000",
16344 => "000010011",
16345 => "000011000",
16346 => "000011101",
16347 => "000101110",
16348 => "000110100",
16349 => "000011101",
16350 => "000110001",
16351 => "001000001",
16352 => "000101111",
16353 => "000110100",
16354 => "001001101",
16355 => "000111010",
16356 => "000100010",
16357 => "001001000",
16358 => "001010110",
16359 => "000110111",
16360 => "001000101",
16361 => "001010000",
16362 => "001011100",
16363 => "001011111",
16364 => "001011011",
16365 => "001010111",
16366 => "001010111",
16367 => "001011001",
16368 => "001010111",
16369 => "001010110",
16370 => "001011000",
16371 => "001010110",
16372 => "001010111",
16373 => "001010001",
16374 => "001010001",
16375 => "001010010",
16376 => "001010110",
16377 => "001001101",
16378 => "001001010",
16379 => "001001001",
16380 => "001001001",
16381 => "001010010",
16382 => "001000111",
16383 => "001001011"
  );

  signal STREAM_0     : std_logic_vector(14 downto 0);
  signal STREAM_0_STB : std_logic;
  signal STREAM_0_ACK : std_logic;

  component RAMARRAY is
    generic(
        DEPTH : integer;
        WIDTH : integer
    );
    port(
        CLK             : in  std_logic;
        RST             : in  std_logic;
        ADDRESS_IN      : in  std_logic_vector;
        ADDRESS_IN_STB  : in  std_logic;
        ADDRESS_IN_ACK  : out std_logic;
        DATA_IN         : in  std_logic_vector;
        DATA_IN_STB     : in  std_logic;
        DATA_IN_ACK     : out std_logic;
        ADDRESS_OUT     : in  std_logic_vector;
        ADDRESS_OUT_STB : in  std_logic;
        ADDRESS_OUT_ACK : out std_logic;
        DATA_OUT        : out std_logic_vector;
        DATA_OUT_STB    : out std_logic;
        DATA_OUT_ACK    : in  std_logic
    );
  end component RAMARRAY;

  signal STREAM_6     : std_logic_vector(12 downto 0);
  signal STREAM_6_STB : std_logic;
  signal STREAM_6_ACK : std_logic;

  signal STREAM_3       : std_logic_vector(12 downto 0);
  signal STREAM_3_STB   : std_logic;
  signal STREAM_3_ACK   : std_logic;
  signal STREAM_4       : std_logic_vector(12 downto 0);
  signal STREAM_4_STB   : std_logic;
  signal STREAM_4_ACK   : std_logic;
  signal STREAM_5       : std_logic_vector(12 downto 0);
  signal STREAM_5_STB   : std_logic;
  signal STREAM_5_ACK   : std_logic;
  signal STREAM_2       : std_logic_vector(12 downto 0);
  signal STREAM_2_STB   : std_logic;
  signal STREAM_2_ACK   : std_logic;
  constant OP_IMM_7 : std_logic_vector(3 downto 0) := "0000";
  constant OP_MOVE_7 : std_logic_vector(3 downto 0) := "0001";
  constant OP_GT_7 : std_logic_vector(3 downto 0) := "0010";
  constant OP_EQ_7 : std_logic_vector(3 downto 0) := "0011";
  constant OP_JMPF_7 : std_logic_vector(3 downto 0) := "0100";
  constant OP_JMP_7 : std_logic_vector(3 downto 0) := "0101";
  constant OP_ADD_7 : std_logic_vector(3 downto 0) := "0110";
  constant OP_GE_7 : std_logic_vector(3 downto 0) := "0111";
  constant OP_SUB_7 : std_logic_vector(3 downto 0) := "1000";
  constant OP_SR_7 : std_logic_vector(3 downto 0) := "1001";
  constant OP_READ_1_7 : std_logic_vector(3 downto 0) := "1010";
  constant OP_READ_6_7 : std_logic_vector(3 downto 0) := "1011";
  constant OP_WRITE_3_7 : std_logic_vector(3 downto 0) := "1100";
  constant OP_WRITE_4_7 : std_logic_vector(3 downto 0) := "1101";
  constant OP_WRITE_5_7 : std_logic_vector(3 downto 0) := "1110";
  constant OP_WRITE_2_7 : std_logic_vector(3 downto 0) := "1111";
  type PROCESS_7_STATE_TYPE is (STALL, EXECUTE, READ_STREAM_1, ACK_STREAM_1, READ_STREAM_6, ACK_STREAM_6, WRITE_STREAM_3, WRITE_STREAM_4, WRITE_STREAM_5, WRITE_STREAM_2);
  type INSTRUCTIONS_TYPE_7  is array (0 to 515) of std_logic_vector(20 downto 0);
  type REGISTERS_TYPE_7     is array (0 to 15) of std_logic_vector(12 downto 0);
  signal STATE_7        : PROCESS_7_STATE_TYPE;
  signal REGISTERS_7    : REGISTERS_TYPE_7;
  signal PC_7           : unsigned(9 downto 0);
  signal OPERATION_7    : std_logic_vector(3 downto 0);
  signal SRCA_7         : std_logic_vector(3 downto 0);
  signal SRCB_7         : std_logic_vector(3 downto 0);
  signal IMMEDIATE_7    : std_logic_vector(12 downto 0);
  signal ZERO_7         : std_logic;
  signal A_7            : std_logic_vector(12 downto 0);
  signal B_7            : std_logic_vector(12 downto 0);
  signal QUOTIENT_7     : std_logic_vector(12 downto 0);
  signal SHIFTER_7      : std_logic_vector(12 downto 0);
  signal REMAINDER_7    : std_logic_vector(12 downto 0);
  signal COUNT_7        : integer range 0 to 13;
  signal SIGN_7         : std_logic;
  signal INSTRUCTIONS_7 : INSTRUCTIONS_TYPE_7 := (
0 => OP_IMM_7 & "0001" & "0000000000000", -- file: ./example_5_edge_detect.py line: 41
1 => OP_IMM_7 & "0010" & "0000000000000", -- file: ./example_5_edge_detect.py line: 43
2 => OP_IMM_7 & "0011" & "0000000000000", -- file: ./example_5_edge_detect.py line: 42
3 => OP_IMM_7 & "0100" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 193
4 => OP_IMM_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
5 => OP_MOVE_7 & "0001" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
6 => OP_IMM_7 & "0101" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
7 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
8 => OP_GT_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
9 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
10 => OP_EQ_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 150
11 => OP_JMPF_7 & "0101" & "0000000001110", -- file: None line: None
12 => OP_JMP_7 & "0000" & "0000000011001", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 63
13 => OP_JMP_7 & "0000" & "0000000001110", -- file: None line: None
14 => OP_IMM_7 & "0101" & "0000100000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
15 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
16 => OP_ADD_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 162
17 => OP_WRITE_3_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
18 => OP_IMM_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
19 => OP_WRITE_4_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
20 => OP_MOVE_7 & "0101" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
21 => OP_IMM_7 & "0110" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
22 => OP_ADD_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
23 => OP_MOVE_7 & "0001" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
24 => OP_JMP_7 & "0000" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 64
25 => OP_IMM_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
26 => OP_MOVE_7 & "0001" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
27 => OP_IMM_7 & "0101" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
28 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
29 => OP_GT_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
30 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
31 => OP_EQ_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 150
32 => OP_JMPF_7 & "0101" & "0000000100011", -- file: None line: None
33 => OP_JMP_7 & "0000" & "0000000101111", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 63
34 => OP_JMP_7 & "0000" & "0000000100011", -- file: None line: None
35 => OP_READ_1_7 & "0010" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 357
36 => OP_IMM_7 & "0101" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
37 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
38 => OP_ADD_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 162
39 => OP_WRITE_3_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
40 => OP_MOVE_7 & "0101" & "0000000000010", -- file: ./example_5_edge_detect.py line: 43
41 => OP_WRITE_4_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
42 => OP_MOVE_7 & "0101" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
43 => OP_IMM_7 & "0110" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
44 => OP_ADD_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
45 => OP_MOVE_7 & "0001" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
46 => OP_JMP_7 & "0000" & "0000000011011", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 64
47 => OP_IMM_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
48 => OP_MOVE_7 & "0001" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
49 => OP_IMM_7 & "0101" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
50 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
51 => OP_GT_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
52 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
53 => OP_EQ_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 150
54 => OP_JMPF_7 & "0101" & "0000000111001", -- file: None line: None
55 => OP_JMP_7 & "0000" & "0000001000011", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 63
56 => OP_JMP_7 & "0000" & "0000000111001", -- file: None line: None
57 => OP_READ_1_7 & "0010" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 357
58 => OP_MOVE_7 & "0101" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
59 => OP_WRITE_3_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
60 => OP_MOVE_7 & "0101" & "0000000000010", -- file: ./example_5_edge_detect.py line: 43
61 => OP_WRITE_4_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
62 => OP_MOVE_7 & "0101" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
63 => OP_IMM_7 & "0110" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
64 => OP_ADD_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
65 => OP_MOVE_7 & "0001" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
66 => OP_JMP_7 & "0000" & "0000000110001", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 64
67 => OP_IMM_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
68 => OP_MOVE_7 & "0011" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
69 => OP_IMM_7 & "0101" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
70 => OP_MOVE_7 & "0110" & "0000000000011", -- file: ./example_5_edge_detect.py line: 42
71 => OP_GT_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
72 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
73 => OP_EQ_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 150
74 => OP_JMPF_7 & "0101" & "0000001001101", -- file: None line: None
75 => OP_JMP_7 & "0000" & "0001000000010", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 63
76 => OP_JMP_7 & "0000" & "0000001001101", -- file: None line: None
77 => OP_IMM_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
78 => OP_MOVE_7 & "0001" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
79 => OP_IMM_7 & "0101" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
80 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
81 => OP_GT_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
82 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
83 => OP_EQ_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 150
84 => OP_JMPF_7 & "0101" & "0000001010111", -- file: None line: None
85 => OP_JMP_7 & "0000" & "0000110100111", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 63
86 => OP_JMP_7 & "0000" & "0000001010111", -- file: None line: None
87 => OP_IMM_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
88 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
89 => OP_GT_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
90 => OP_JMPF_7 & "0101" & "0000001011111", -- file: None line: None
91 => OP_IMM_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
92 => OP_MOVE_7 & "0000" & "0000000000101", -- file: ./example_5_edge_detect.py line: 36
93 => OP_JMP_7 & "0000" & "0000001110010", -- file: ./example_5_edge_detect.py line: 36
94 => OP_JMP_7 & "0000" & "0000001011111", -- file: None line: None
95 => OP_MOVE_7 & "0101" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
96 => OP_IMM_7 & "0110" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
97 => OP_GE_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 156
98 => OP_JMPF_7 & "0101" & "0000001100111", -- file: None line: None
99 => OP_IMM_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
100 => OP_MOVE_7 & "0000" & "0000000000101", -- file: ./example_5_edge_detect.py line: 37
101 => OP_JMP_7 & "0000" & "0000001110010", -- file: ./example_5_edge_detect.py line: 37
102 => OP_JMP_7 & "0000" & "0000001100111", -- file: None line: None
103 => OP_MOVE_7 & "0101" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
104 => OP_IMM_7 & "0110" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
105 => OP_ADD_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
106 => OP_WRITE_5_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
107 => OP_READ_6_7 & "0100" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 357
108 => OP_MOVE_7 & "0101" & "0000000000100", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 193
109 => OP_MOVE_7 & "0000" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
110 => OP_JMP_7 & "0000" & "0000001101111", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
111 => OP_MOVE_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
112 => OP_MOVE_7 & "0000" & "0000000000101", -- file: ./example_5_edge_detect.py line: 38
113 => OP_JMP_7 & "0000" & "0000001110010", -- file: ./example_5_edge_detect.py line: 38
114 => OP_MOVE_7 & "0101" & "0000000000000", -- file: ./example_5_edge_detect.py line: 38
115 => OP_MOVE_7 & "0010" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
116 => OP_MOVE_7 & "0101" & "0000000000010", -- file: ./example_5_edge_detect.py line: 43
117 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
118 => OP_MOVE_7 & "0111" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
119 => OP_IMM_7 & "1000" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
120 => OP_SUB_7 & "0111" & "0000000001000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 132
121 => OP_GT_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
122 => OP_JMPF_7 & "0110" & "0000001111111", -- file: None line: None
123 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
124 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 36
125 => OP_JMP_7 & "0000" & "0000010010110", -- file: ./example_5_edge_detect.py line: 36
126 => OP_JMP_7 & "0000" & "0000001111111", -- file: None line: None
127 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
128 => OP_IMM_7 & "0111" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
129 => OP_SUB_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 132
130 => OP_IMM_7 & "0111" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
131 => OP_GE_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 156
132 => OP_JMPF_7 & "0110" & "0000010001001", -- file: None line: None
133 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
134 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 37
135 => OP_JMP_7 & "0000" & "0000010010110", -- file: ./example_5_edge_detect.py line: 37
136 => OP_JMP_7 & "0000" & "0000010001001", -- file: None line: None
137 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
138 => OP_IMM_7 & "0111" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
139 => OP_SUB_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 132
140 => OP_IMM_7 & "0111" & "0000100000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
141 => OP_ADD_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
142 => OP_WRITE_5_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
143 => OP_READ_6_7 & "0100" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 357
144 => OP_MOVE_7 & "0110" & "0000000000100", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 193
145 => OP_MOVE_7 & "0000" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
146 => OP_JMP_7 & "0000" & "0000010010011", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
147 => OP_MOVE_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
148 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 38
149 => OP_JMP_7 & "0000" & "0000010010110", -- file: ./example_5_edge_detect.py line: 38
150 => OP_MOVE_7 & "0110" & "0000000000000", -- file: ./example_5_edge_detect.py line: 38
151 => OP_IMM_7 & "0111" & "0000000000011", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
152 => OP_SR_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 146
153 => OP_SUB_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 132
154 => OP_MOVE_7 & "0010" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
155 => OP_MOVE_7 & "0101" & "0000000000010", -- file: ./example_5_edge_detect.py line: 43
156 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
157 => OP_MOVE_7 & "0111" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
158 => OP_IMM_7 & "1000" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
159 => OP_SUB_7 & "0111" & "0000000001000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 132
160 => OP_GT_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
161 => OP_JMPF_7 & "0110" & "0000010100110", -- file: None line: None
162 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
163 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 36
164 => OP_JMP_7 & "0000" & "0000010111101", -- file: ./example_5_edge_detect.py line: 36
165 => OP_JMP_7 & "0000" & "0000010100110", -- file: None line: None
166 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
167 => OP_IMM_7 & "0111" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
168 => OP_SUB_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 132
169 => OP_IMM_7 & "0111" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
170 => OP_GE_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 156
171 => OP_JMPF_7 & "0110" & "0000010110000", -- file: None line: None
172 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
173 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 37
174 => OP_JMP_7 & "0000" & "0000010111101", -- file: ./example_5_edge_detect.py line: 37
175 => OP_JMP_7 & "0000" & "0000010110000", -- file: None line: None
176 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
177 => OP_IMM_7 & "0111" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
178 => OP_SUB_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 132
179 => OP_IMM_7 & "0111" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
180 => OP_ADD_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
181 => OP_WRITE_5_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
182 => OP_READ_6_7 & "0100" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 357
183 => OP_MOVE_7 & "0110" & "0000000000100", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 193
184 => OP_MOVE_7 & "0000" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
185 => OP_JMP_7 & "0000" & "0000010111010", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
186 => OP_MOVE_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
187 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 38
188 => OP_JMP_7 & "0000" & "0000010111101", -- file: ./example_5_edge_detect.py line: 38
189 => OP_MOVE_7 & "0110" & "0000000000000", -- file: ./example_5_edge_detect.py line: 38
190 => OP_IMM_7 & "0111" & "0000000000011", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
191 => OP_SR_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 146
192 => OP_SUB_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 132
193 => OP_MOVE_7 & "0010" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
194 => OP_MOVE_7 & "0101" & "0000000000010", -- file: ./example_5_edge_detect.py line: 43
195 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
196 => OP_MOVE_7 & "0111" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
197 => OP_IMM_7 & "1000" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
198 => OP_SUB_7 & "0111" & "0000000001000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 132
199 => OP_GT_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
200 => OP_JMPF_7 & "0110" & "0000011001101", -- file: None line: None
201 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
202 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 36
203 => OP_JMP_7 & "0000" & "0000011100100", -- file: ./example_5_edge_detect.py line: 36
204 => OP_JMP_7 & "0000" & "0000011001101", -- file: None line: None
205 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
206 => OP_IMM_7 & "0111" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
207 => OP_SUB_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 132
208 => OP_IMM_7 & "0111" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
209 => OP_GE_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 156
210 => OP_JMPF_7 & "0110" & "0000011010111", -- file: None line: None
211 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
212 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 37
213 => OP_JMP_7 & "0000" & "0000011100100", -- file: ./example_5_edge_detect.py line: 37
214 => OP_JMP_7 & "0000" & "0000011010111", -- file: None line: None
215 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
216 => OP_IMM_7 & "0111" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
217 => OP_SUB_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 132
218 => OP_IMM_7 & "0111" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
219 => OP_ADD_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
220 => OP_WRITE_5_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
221 => OP_READ_6_7 & "0100" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 357
222 => OP_MOVE_7 & "0110" & "0000000000100", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 193
223 => OP_MOVE_7 & "0000" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
224 => OP_JMP_7 & "0000" & "0000011100001", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
225 => OP_MOVE_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
226 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 38
227 => OP_JMP_7 & "0000" & "0000011100100", -- file: ./example_5_edge_detect.py line: 38
228 => OP_MOVE_7 & "0110" & "0000000000000", -- file: ./example_5_edge_detect.py line: 38
229 => OP_IMM_7 & "0111" & "0000000000011", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
230 => OP_SR_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 146
231 => OP_SUB_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 132
232 => OP_MOVE_7 & "0010" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
233 => OP_MOVE_7 & "0101" & "0000000000010", -- file: ./example_5_edge_detect.py line: 43
234 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
235 => OP_MOVE_7 & "0111" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
236 => OP_GT_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
237 => OP_JMPF_7 & "0110" & "0000011110010", -- file: None line: None
238 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
239 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 36
240 => OP_JMP_7 & "0000" & "0000100000101", -- file: ./example_5_edge_detect.py line: 36
241 => OP_JMP_7 & "0000" & "0000011110010", -- file: None line: None
242 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
243 => OP_IMM_7 & "0111" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
244 => OP_GE_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 156
245 => OP_JMPF_7 & "0110" & "0000011111010", -- file: None line: None
246 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
247 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 37
248 => OP_JMP_7 & "0000" & "0000100000101", -- file: ./example_5_edge_detect.py line: 37
249 => OP_JMP_7 & "0000" & "0000011111010", -- file: None line: None
250 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
251 => OP_IMM_7 & "0111" & "0000100000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
252 => OP_ADD_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
253 => OP_WRITE_5_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
254 => OP_READ_6_7 & "0100" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 357
255 => OP_MOVE_7 & "0110" & "0000000000100", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 193
256 => OP_MOVE_7 & "0000" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
257 => OP_JMP_7 & "0000" & "0000100000010", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
258 => OP_MOVE_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
259 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 38
260 => OP_JMP_7 & "0000" & "0000100000101", -- file: ./example_5_edge_detect.py line: 38
261 => OP_MOVE_7 & "0110" & "0000000000000", -- file: ./example_5_edge_detect.py line: 38
262 => OP_IMM_7 & "0111" & "0000000000011", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
263 => OP_SR_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 146
264 => OP_SUB_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 132
265 => OP_MOVE_7 & "0010" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
266 => OP_MOVE_7 & "0101" & "0000000000010", -- file: ./example_5_edge_detect.py line: 43
267 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
268 => OP_MOVE_7 & "0111" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
269 => OP_GT_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
270 => OP_JMPF_7 & "0110" & "0000100010011", -- file: None line: None
271 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
272 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 36
273 => OP_JMP_7 & "0000" & "0000100100110", -- file: ./example_5_edge_detect.py line: 36
274 => OP_JMP_7 & "0000" & "0000100010011", -- file: None line: None
275 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
276 => OP_IMM_7 & "0111" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
277 => OP_GE_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 156
278 => OP_JMPF_7 & "0110" & "0000100011011", -- file: None line: None
279 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
280 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 37
281 => OP_JMP_7 & "0000" & "0000100100110", -- file: ./example_5_edge_detect.py line: 37
282 => OP_JMP_7 & "0000" & "0000100011011", -- file: None line: None
283 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
284 => OP_IMM_7 & "0111" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
285 => OP_ADD_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
286 => OP_WRITE_5_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
287 => OP_READ_6_7 & "0100" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 357
288 => OP_MOVE_7 & "0110" & "0000000000100", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 193
289 => OP_MOVE_7 & "0000" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
290 => OP_JMP_7 & "0000" & "0000100100011", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
291 => OP_MOVE_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
292 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 38
293 => OP_JMP_7 & "0000" & "0000100100110", -- file: ./example_5_edge_detect.py line: 38
294 => OP_MOVE_7 & "0110" & "0000000000000", -- file: ./example_5_edge_detect.py line: 38
295 => OP_IMM_7 & "0111" & "0000000000011", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
296 => OP_SR_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 146
297 => OP_SUB_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 132
298 => OP_MOVE_7 & "0010" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
299 => OP_MOVE_7 & "0101" & "0000000000010", -- file: ./example_5_edge_detect.py line: 43
300 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
301 => OP_MOVE_7 & "0111" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
302 => OP_IMM_7 & "1000" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
303 => OP_ADD_7 & "0111" & "0000000001000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
304 => OP_GT_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
305 => OP_JMPF_7 & "0110" & "0000100110110", -- file: None line: None
306 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
307 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 36
308 => OP_JMP_7 & "0000" & "0000101001101", -- file: ./example_5_edge_detect.py line: 36
309 => OP_JMP_7 & "0000" & "0000100110110", -- file: None line: None
310 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
311 => OP_IMM_7 & "0111" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
312 => OP_ADD_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
313 => OP_IMM_7 & "0111" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
314 => OP_GE_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 156
315 => OP_JMPF_7 & "0110" & "0000101000000", -- file: None line: None
316 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
317 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 37
318 => OP_JMP_7 & "0000" & "0000101001101", -- file: ./example_5_edge_detect.py line: 37
319 => OP_JMP_7 & "0000" & "0000101000000", -- file: None line: None
320 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
321 => OP_IMM_7 & "0111" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
322 => OP_ADD_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
323 => OP_IMM_7 & "0111" & "0000100000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
324 => OP_ADD_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
325 => OP_WRITE_5_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
326 => OP_READ_6_7 & "0100" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 357
327 => OP_MOVE_7 & "0110" & "0000000000100", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 193
328 => OP_MOVE_7 & "0000" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
329 => OP_JMP_7 & "0000" & "0000101001010", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
330 => OP_MOVE_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
331 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 38
332 => OP_JMP_7 & "0000" & "0000101001101", -- file: ./example_5_edge_detect.py line: 38
333 => OP_MOVE_7 & "0110" & "0000000000000", -- file: ./example_5_edge_detect.py line: 38
334 => OP_IMM_7 & "0111" & "0000000000011", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
335 => OP_SR_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 146
336 => OP_SUB_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 132
337 => OP_MOVE_7 & "0010" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
338 => OP_MOVE_7 & "0101" & "0000000000010", -- file: ./example_5_edge_detect.py line: 43
339 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
340 => OP_MOVE_7 & "0111" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
341 => OP_IMM_7 & "1000" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
342 => OP_ADD_7 & "0111" & "0000000001000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
343 => OP_GT_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
344 => OP_JMPF_7 & "0110" & "0000101011101", -- file: None line: None
345 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
346 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 36
347 => OP_JMP_7 & "0000" & "0000101110100", -- file: ./example_5_edge_detect.py line: 36
348 => OP_JMP_7 & "0000" & "0000101011101", -- file: None line: None
349 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
350 => OP_IMM_7 & "0111" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
351 => OP_ADD_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
352 => OP_IMM_7 & "0111" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
353 => OP_GE_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 156
354 => OP_JMPF_7 & "0110" & "0000101100111", -- file: None line: None
355 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
356 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 37
357 => OP_JMP_7 & "0000" & "0000101110100", -- file: ./example_5_edge_detect.py line: 37
358 => OP_JMP_7 & "0000" & "0000101100111", -- file: None line: None
359 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
360 => OP_IMM_7 & "0111" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
361 => OP_ADD_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
362 => OP_IMM_7 & "0111" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
363 => OP_ADD_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
364 => OP_WRITE_5_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
365 => OP_READ_6_7 & "0100" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 357
366 => OP_MOVE_7 & "0110" & "0000000000100", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 193
367 => OP_MOVE_7 & "0000" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
368 => OP_JMP_7 & "0000" & "0000101110001", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
369 => OP_MOVE_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
370 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 38
371 => OP_JMP_7 & "0000" & "0000101110100", -- file: ./example_5_edge_detect.py line: 38
372 => OP_MOVE_7 & "0110" & "0000000000000", -- file: ./example_5_edge_detect.py line: 38
373 => OP_IMM_7 & "0111" & "0000000000011", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
374 => OP_SR_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 146
375 => OP_SUB_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 132
376 => OP_MOVE_7 & "0010" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
377 => OP_MOVE_7 & "0101" & "0000000000010", -- file: ./example_5_edge_detect.py line: 43
378 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
379 => OP_MOVE_7 & "0111" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
380 => OP_IMM_7 & "1000" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
381 => OP_ADD_7 & "0111" & "0000000001000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
382 => OP_GT_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
383 => OP_JMPF_7 & "0110" & "0000110000100", -- file: None line: None
384 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
385 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 36
386 => OP_JMP_7 & "0000" & "0000110011011", -- file: ./example_5_edge_detect.py line: 36
387 => OP_JMP_7 & "0000" & "0000110000100", -- file: None line: None
388 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
389 => OP_IMM_7 & "0111" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
390 => OP_ADD_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
391 => OP_IMM_7 & "0111" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
392 => OP_GE_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 156
393 => OP_JMPF_7 & "0110" & "0000110001110", -- file: None line: None
394 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
395 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 37
396 => OP_JMP_7 & "0000" & "0000110011011", -- file: ./example_5_edge_detect.py line: 37
397 => OP_JMP_7 & "0000" & "0000110001110", -- file: None line: None
398 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
399 => OP_IMM_7 & "0111" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
400 => OP_ADD_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
401 => OP_IMM_7 & "0111" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
402 => OP_ADD_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
403 => OP_WRITE_5_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
404 => OP_READ_6_7 & "0100" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 357
405 => OP_MOVE_7 & "0110" & "0000000000100", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 193
406 => OP_MOVE_7 & "0000" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
407 => OP_JMP_7 & "0000" & "0000110011000", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
408 => OP_MOVE_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
409 => OP_MOVE_7 & "0000" & "0000000000110", -- file: ./example_5_edge_detect.py line: 38
410 => OP_JMP_7 & "0000" & "0000110011011", -- file: ./example_5_edge_detect.py line: 38
411 => OP_MOVE_7 & "0110" & "0000000000000", -- file: ./example_5_edge_detect.py line: 38
412 => OP_IMM_7 & "0111" & "0000000000011", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
413 => OP_SR_7 & "0110" & "0000000000111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 146
414 => OP_SUB_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 132
415 => OP_MOVE_7 & "0010" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
416 => OP_MOVE_7 & "0101" & "0000000000010", -- file: ./example_5_edge_detect.py line: 43
417 => OP_WRITE_2_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
418 => OP_MOVE_7 & "0101" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
419 => OP_IMM_7 & "0110" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
420 => OP_ADD_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
421 => OP_MOVE_7 & "0001" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
422 => OP_JMP_7 & "0000" & "0000001001111", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 64
423 => OP_IMM_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
424 => OP_MOVE_7 & "0001" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
425 => OP_IMM_7 & "0101" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
426 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
427 => OP_GT_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
428 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
429 => OP_EQ_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 150
430 => OP_JMPF_7 & "0101" & "0000110110001", -- file: None line: None
431 => OP_JMP_7 & "0000" & "0000111000100", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 63
432 => OP_JMP_7 & "0000" & "0000110110001", -- file: None line: None
433 => OP_IMM_7 & "0101" & "0000100000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
434 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
435 => OP_ADD_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 162
436 => OP_WRITE_3_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
437 => OP_IMM_7 & "0101" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
438 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
439 => OP_ADD_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 162
440 => OP_WRITE_5_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
441 => OP_READ_6_7 & "0100" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 357
442 => OP_MOVE_7 & "0101" & "0000000000100", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 193
443 => OP_MOVE_7 & "0000" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
444 => OP_JMP_7 & "0000" & "0000110111101", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
445 => OP_MOVE_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
446 => OP_WRITE_4_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
447 => OP_MOVE_7 & "0101" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
448 => OP_IMM_7 & "0110" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
449 => OP_ADD_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
450 => OP_MOVE_7 & "0001" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
451 => OP_JMP_7 & "0000" & "0000110101001", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 64
452 => OP_IMM_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
453 => OP_MOVE_7 & "0001" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
454 => OP_IMM_7 & "0101" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
455 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
456 => OP_GT_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
457 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
458 => OP_EQ_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 150
459 => OP_JMPF_7 & "0101" & "0000111001110", -- file: None line: None
460 => OP_JMP_7 & "0000" & "0000111011111", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 63
461 => OP_JMP_7 & "0000" & "0000111001110", -- file: None line: None
462 => OP_IMM_7 & "0101" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
463 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
464 => OP_ADD_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 162
465 => OP_WRITE_3_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
466 => OP_MOVE_7 & "0101" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
467 => OP_WRITE_5_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
468 => OP_READ_6_7 & "0100" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 357
469 => OP_MOVE_7 & "0101" & "0000000000100", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 193
470 => OP_MOVE_7 & "0000" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
471 => OP_JMP_7 & "0000" & "0000111011000", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
472 => OP_MOVE_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 204
473 => OP_WRITE_4_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
474 => OP_MOVE_7 & "0101" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
475 => OP_IMM_7 & "0110" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
476 => OP_ADD_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
477 => OP_MOVE_7 & "0001" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
478 => OP_JMP_7 & "0000" & "0000111000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 64
479 => OP_IMM_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
480 => OP_MOVE_7 & "0001" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
481 => OP_IMM_7 & "0101" & "0000010000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
482 => OP_MOVE_7 & "0110" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
483 => OP_GT_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
484 => OP_IMM_7 & "0110" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
485 => OP_EQ_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 150
486 => OP_JMPF_7 & "0101" & "0000111101001", -- file: None line: None
487 => OP_JMP_7 & "0000" & "0000111111101", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 63
488 => OP_JMP_7 & "0000" & "0000111101001", -- file: None line: None
489 => OP_IMM_7 & "0101" & "0000001111111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
490 => OP_MOVE_7 & "0110" & "0000000000011", -- file: ./example_5_edge_detect.py line: 42
491 => OP_GT_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 158
492 => OP_JMPF_7 & "0101" & "0000111101111", -- file: None line: None
493 => OP_READ_1_7 & "0010" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 357
494 => OP_JMP_7 & "0000" & "0000111110100", -- file: None line: None
495 => OP_IMM_7 & "0101" & "1111111111111", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
496 => OP_JMPF_7 & "0101" & "0000111110100", -- file: None line: None
497 => OP_IMM_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
498 => OP_MOVE_7 & "0010" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
499 => OP_JMP_7 & "0000" & "0000111110100", -- file: None line: None
500 => OP_MOVE_7 & "0101" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
501 => OP_WRITE_3_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
502 => OP_MOVE_7 & "0101" & "0000000000010", -- file: ./example_5_edge_detect.py line: 43
503 => OP_WRITE_4_7 & "0101" & "0000000000000", -- file: /usr/local/lib/python2.6/dist-packages/chips/streams.py line: 715
504 => OP_MOVE_7 & "0101" & "0000000000001", -- file: ./example_5_edge_detect.py line: 41
505 => OP_IMM_7 & "0110" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
506 => OP_ADD_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
507 => OP_MOVE_7 & "0001" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
508 => OP_JMP_7 & "0000" & "0000111100001", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 64
509 => OP_MOVE_7 & "0101" & "0000000000011", -- file: ./example_5_edge_detect.py line: 42
510 => OP_IMM_7 & "0110" & "0000000000001", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 114
511 => OP_ADD_7 & "0101" & "0000000000110", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 130
512 => OP_MOVE_7 & "0011" & "0000000000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/instruction.py line: 375
513 => OP_JMP_7 & "0000" & "0000001000101", -- file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py line: 64
514 => OP_JMP_7 & "0000" & "0001000000010", -- file: None line: None
515 => OP_JMP_7 & "0000" & "0000000000000"); -- file: None line: None
  signal MOD_DIV_7      : std_logic;

begin

  process
  begin
    wait until rising_edge(CLK);
    TIMER_1us <= '0';
    TIMER_10us <= '0';
    TIMER_100us <= '0';
    TIMER_1ms <= '0';
    if TIMER_1us_COUNT = 0 then
       TIMER_1us_COUNT <= TIMER_1us_MAX;
       TIMER_1us <= '1';
       if TIMER_10us_COUNT = 0 then
         TIMER_10us_COUNT <= TIMER_10us_MAX;
         TIMER_10us <= '1';
         if TIMER_100us_COUNT = 0 then
           TIMER_100us_COUNT <= TIMER_100us_MAX;
           TIMER_100us <= '1';
           if TIMER_1ms_COUNT = 0 then
             TIMER_1ms_COUNT <= TIMER_1ms_MAX;
             TIMER_1ms <= '1';
           else
             TIMER_1ms_COUNT <= TIMER_1ms_COUNT - 1;
           end if;
         else
           TIMER_100us_COUNT <= TIMER_100us_COUNT - 1;
         end if;
       else
         TIMER_10us_COUNT <= TIMER_10us_COUNT - 1;
       end if;
    else
       TIMER_1us_COUNT <= TIMER_1us_COUNT - 1;
    end if;
    if RST = '1' then
       TIMER_1us_COUNT <= TIMER_1us_MAX;
       TIMER_1us <= '0';
       TIMER_10us_COUNT <= TIMER_10us_MAX;
       TIMER_10us <= '0';
       TIMER_100us_COUNT <= TIMER_100us_MAX;
       TIMER_100us <= '0';
       TIMER_1ms_COUNT <= TIMER_1ms_MAX;
       TIMER_1ms <= '0';
    end if;
  end process;

  --internal clock generator
  process
  begin
    while True loop
      CLK <= '0';
      wait for 5 ns;
      CLK <= '1';
      wait for 5 ns;
    end loop;
    wait;
  end process;

  --internal reset generator
  process
  begin
    RST <= '1';
    wait for 20 ns;
    RST <= '0';
    wait;
  end process;

  --file: ./example_5_edge_detect.py, line: 156
  --OutPort(2, 13)
  process
    file OUTFILE : text open write_mode is "resp_2.txt";
    variable OUTLINE : LINE;
    variable VALUE : integer;
  begin
    wait until rising_edge(CLK);
    STREAM_2_ACK <= '0';
    if STREAM_2_STB = '1' then
      STREAM_2_ACK <= '1';
    end if;    if STREAM_2_STB = '1' and STREAM_2_ACK = '1' then
      VALUE := to_integer(signed(STREAM_2));
      write(OUTLINE, VALUE);
      writeline(OUTFILE, OUTLINE);
    end if;  end process;

  --file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py, line: 59
  --STREAM 1 Lookup()
  process
  begin
    wait until rising_edge(CLK);
    case STATE_1 is
      when UNARY_INPUT =>
        if STREAM_0_STB = '1' then
          STREAM_0_ACK <= '1';
          STREAM_1_STB <= '1';
          STREAM_1 <= LOOKUP_1(to_integer(unsigned(STREAM_0)));
          STATE_1 <= UNARY_OUTPUT;
        end if;
      when UNARY_OUTPUT =>
        STREAM_0_ACK <= '0';
        if STREAM_1_ACK = '1' then
           STREAM_1_STB <= '0';
           STATE_1 <= UNARY_INPUT;
        end if;
     end case;
     if RST = '1' then
       STREAM_1_STB <= '0';
       STREAM_0_ACK <= '0';
       STATE_1 <= UNARY_INPUT;
     end if;
  end process;

  --file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py, line: 59
  --STREAM 0 Counter(0, 16383, 1, 15)
  process
  begin
    wait until rising_edge(CLK);
    STREAM_0_STB <= '1';
    if STREAM_0_ACK = '1' then
      STREAM_0_STB <= '0';
      STREAM_0 <= STD_RESIZE(ADD(STREAM_0, "000000000000001"), 15);
      if STREAM_0 = "011111111111111" then
        STREAM_0 <= "000000000000000";
      end if;
    end if;
    if RST = '1' then
      STREAM_0_STB <= '0';
      STREAM_0 <= "000000000000000";
    end if;
  end process;

  --file: /usr/local/lib/python2.6/dist-packages/chips/__init__.py, line: 194
  --STREAM 6 Array()
    RAMARRAY_6 : RAMARRAY generic map(
      DEPTH => 384,
      WIDTH => 13
    )
    port map(
      CLK             => CLK,
      RST             => RST,
      ADDRESS_IN      => STREAM_3,
      ADDRESS_IN_STB  => STREAM_3_STB,
      ADDRESS_IN_ACK  => STREAM_3_ACK,
      DATA_IN         => STREAM_4,
      DATA_IN_STB     => STREAM_4_STB,
      DATA_IN_ACK     => STREAM_4_ACK,
      ADDRESS_OUT     => STREAM_5,
      ADDRESS_OUT_STB => STREAM_5_STB,
      ADDRESS_OUT_ACK => STREAM_5_ACK,
      DATA_OUT        => STREAM_6,
      DATA_OUT_STB    => STREAM_6_STB,
      DATA_OUT_ACK    => STREAM_6_ACK
    );

  -- process
  process
    variable INSTRUCTION : std_logic_vector(20 downto 0);
  begin
    wait until rising_edge(CLK);
    INSTRUCTION := INSTRUCTIONS_7(to_integer(PC_7));
    OPERATION_7 <= INSTRUCTION(20 downto 17);
    SRCA_7      <= INSTRUCTION(16 downto 13);
    SRCB_7      <= INSTRUCTION(3 downto 0);
    IMMEDIATE_7 <= INSTRUCTION(12 downto 0);
  end process;

  process
    variable REGA         : std_logic_vector(12 downto 0);
    variable REGB         : std_logic_vector(12 downto 0);
    variable DEST         : std_logic_vector(3 downto 0);
    variable RESULT       : std_logic_vector(12 downto 0);
    variable RESULT_DEL   : std_logic_vector(12 downto 0);
    variable REGISTERS_EN : std_logic;
    variable MODULO       : unsigned(12 downto 0);
    variable FLAG_EQ      : std_logic;
    variable FLAG_GT      : std_logic;
    variable FLAG_GE      : std_logic;
  begin
    wait until rising_edge(CLK);
    REGISTERS_EN := '0';
    case STATE_7 is
      when STALL =>
        PC_7 <= PC_7 + 1;
        STATE_7 <= EXECUTE;
      when EXECUTE =>
        REGA := REGISTERS_7(to_integer(unsigned(SRCA_7)));
        REGB := REGISTERS_7(to_integer(unsigned(SRCB_7)));
        DEST := SRCA_7;
        RESULT := REGA;
        PC_7 <= PC_7 + 1;

        --share comparator logic
        if REGA = REGB then
          FLAG_EQ := '1';
        else
          FLAG_EQ := '0';
        end if;

        if signed(REGA) > signed(REGB) then
          FLAG_GT := '1';
        else
          FLAG_GT := '0';
        end if;

        FLAG_GE := FLAG_GT or FLAG_EQ;

        --execute instructions
        case OPERATION_7 is
          when OP_MOVE_7 => 
            RESULT := REGB;
            REGISTERS_EN := '1';
          when OP_ADD_7  => 
            RESULT := STD_RESIZE( ADD(REGA, REGB), 13);
            REGISTERS_EN := '1';
          when OP_SUB_7  => 
            RESULT := STD_RESIZE( SUB(REGA, REGB), 13);
            REGISTERS_EN := '1';
          when OP_SR_7   => 
            RESULT := STD_RESIZE(  SR(REGA, REGB), 13);
            REGISTERS_EN := '1';
          when OP_EQ_7   => 
            RESULT := (others => FLAG_EQ);
            REGISTERS_EN := '1';
          when OP_GT_7   => 
            RESULT := (others => FLAG_GT);
            REGISTERS_EN := '1';
          when OP_GE_7   => 
            RESULT := (others => FLAG_GE);
            REGISTERS_EN := '1';
          when OP_IMM_7  => 
            RESULT := IMMEDIATE_7;
            REGISTERS_EN := '1';
          when OP_JMP_7 =>
            STATE_7 <= STALL;
            PC_7 <= resize(unsigned(IMMEDIATE_7), 10);
          when OP_JMPF_7 =>
            if RESULT_DEL = "0000000000000" then
              STATE_7 <= STALL;
              PC_7 <= resize(unsigned(IMMEDIATE_7), 10);
            end if;

          when OP_WRITE_3_7 =>
            STATE_7 <= WRITE_STREAM_3;
            DEST := SRCA_7;
            PC_7 <= PC_7;
          when OP_WRITE_4_7 =>
            STATE_7 <= WRITE_STREAM_4;
            DEST := SRCA_7;
            PC_7 <= PC_7;
          when OP_WRITE_5_7 =>
            STATE_7 <= WRITE_STREAM_5;
            DEST := SRCA_7;
            PC_7 <= PC_7;
          when OP_WRITE_2_7 =>
            STATE_7 <= WRITE_STREAM_2;
            DEST := SRCA_7;
            PC_7 <= PC_7;
          when OP_READ_1_7 =>
            STATE_7 <= READ_STREAM_1;
            PC_7 <= PC_7;
          when OP_READ_6_7 =>
            STATE_7 <= READ_STREAM_6;
            PC_7 <= PC_7;
          when others => null;
        end case;

        --write back results
        RESULT_DEL := RESULT;

      when READ_STREAM_1 =>
        if STREAM_1_STB = '1' then
          STREAM_1_ACK <= '1';
          REGISTERS_EN := '1';
          RESULT := STD_RESIZE(STREAM_1, 13);
          STATE_7 <= ACK_STREAM_1;
        end if;
      when ACK_STREAM_1 =>
        STREAM_1_ACK <= '0';
        STATE_7 <= EXECUTE;
        PC_7 <= PC_7 + 1;
      when READ_STREAM_6 =>
        if STREAM_6_STB = '1' then
          STREAM_6_ACK <= '1';
          REGISTERS_EN := '1';
          RESULT := STD_RESIZE(STREAM_6, 13);
          STATE_7 <= ACK_STREAM_6;
        end if;
      when ACK_STREAM_6 =>
        STREAM_6_ACK <= '0';
        STATE_7 <= EXECUTE;
        PC_7 <= PC_7 + 1;
      when WRITE_STREAM_3 =>
        STREAM_3_STB <= '1';
        STREAM_3 <= STD_RESIZE(REGA, 13);
        if STREAM_3_ACK = '1' then
          STREAM_3_STB <= '0';
          STATE_7 <= EXECUTE;
          PC_7 <= PC_7 + 1;
        end if;
      when WRITE_STREAM_4 =>
        STREAM_4_STB <= '1';
        STREAM_4 <= STD_RESIZE(REGA, 13);
        if STREAM_4_ACK = '1' then
          STREAM_4_STB <= '0';
          STATE_7 <= EXECUTE;
          PC_7 <= PC_7 + 1;
        end if;
      when WRITE_STREAM_5 =>
        STREAM_5_STB <= '1';
        STREAM_5 <= STD_RESIZE(REGA, 13);
        if STREAM_5_ACK = '1' then
          STREAM_5_STB <= '0';
          STATE_7 <= EXECUTE;
          PC_7 <= PC_7 + 1;
        end if;
      when WRITE_STREAM_2 =>
        STREAM_2_STB <= '1';
        STREAM_2 <= STD_RESIZE(REGA, 13);
        if STREAM_2_ACK = '1' then
          STREAM_2_STB <= '0';
          STATE_7 <= EXECUTE;
          PC_7 <= PC_7 + 1;
        end if;
    end case;

    if RST = '1' then
      STATE_7 <= STALL;
      PC_7 <= "0000000000";
      STREAM_1_ACK <= '0';
      STREAM_6_ACK <= '0';
      STREAM_3_STB <= '0';
      STREAM_4_STB <= '0';
      STREAM_5_STB <= '0';
      STREAM_2_STB <= '0';
    end if;
    if REGISTERS_EN = '1' then
      REGISTERS_7(to_integer(unsigned(DEST))) <= RESULT;
    end if;
  end process;



end architecture RTL;

--+============================================================================+
--|                       **END OF AUTO GENERATED CODE**                       |
--+============================================================================+